-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"f2040000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"8bfc7383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040ba0",
    29 => x"8080fd0b",
    30 => x"a0808bb9",
    31 => x"040ba080",
    32 => x"80fd0402",
    33 => x"c0050d02",
    34 => x"80c40580",
    35 => x"e05c5c80",
    36 => x"7c708405",
    37 => x"5e08715f",
    38 => x"5f587d70",
    39 => x"84055f08",
    40 => x"57805a76",
    41 => x"982a7788",
    42 => x"2b585574",
    43 => x"802e828d",
    44 => x"387c802e",
    45 => x"bf38805d",
    46 => x"7480e42e",
    47 => x"81af3874",
    48 => x"80e42680",
    49 => x"e8387480",
    50 => x"e32e80c1",
    51 => x"38a551a0",
    52 => x"8086a22d",
    53 => x"7451a080",
    54 => x"86a22d82",
    55 => x"1858811a",
    56 => x"5a837a25",
    57 => x"ffbd3874",
    58 => x"ffb0387e",
    59 => x"800c0280",
    60 => x"c0050d04",
    61 => x"74a52e09",
    62 => x"81069a38",
    63 => x"810b811b",
    64 => x"5b5d837a",
    65 => x"25ff9c38",
    66 => x"a08081e7",
    67 => x"047b841d",
    68 => x"7108575d",
    69 => x"547451a0",
    70 => x"8086a22d",
    71 => x"8118811b",
    72 => x"5b58837a",
    73 => x"25fefc38",
    74 => x"a08081e7",
    75 => x"047480f3",
    76 => x"2e098106",
    77 => x"ff97387b",
    78 => x"841d7108",
    79 => x"70545d5d",
    80 => x"53a08088",
    81 => x"be2d800b",
    82 => x"ff115452",
    83 => x"807225ff",
    84 => x"8d387a70",
    85 => x"81055c33",
    86 => x"705255a0",
    87 => x"8086a22d",
    88 => x"811873ff",
    89 => x"15555358",
    90 => x"a08082cc",
    91 => x"047b841d",
    92 => x"71087f5c",
    93 => x"555d5287",
    94 => x"56729c2a",
    95 => x"73842b54",
    96 => x"5271802e",
    97 => x"83388159",
    98 => x"b7125471",
    99 => x"89248438",
   100 => x"b0125478",
   101 => x"9438ff16",
   102 => x"56758025",
   103 => x"dc38800b",
   104 => x"ff115452",
   105 => x"a08082cc",
   106 => x"047351a0",
   107 => x"8086a22d",
   108 => x"ff165675",
   109 => x"8025c238",
   110 => x"a080839e",
   111 => x"0477800c",
   112 => x"0280c005",
   113 => x"0d04830b",
   114 => x"85ffc481",
   115 => x"34fc0b85",
   116 => x"ffc08134",
   117 => x"0402f405",
   118 => x"0dfea080",
   119 => x"0b86ffe2",
   120 => x"8023800b",
   121 => x"86ffe282",
   122 => x"23800b86",
   123 => x"ffe28423",
   124 => x"800b86ff",
   125 => x"e2882380",
   126 => x"0b86ffe2",
   127 => x"8a2381a0",
   128 => x"705353a0",
   129 => x"bf518072",
   130 => x"70840554",
   131 => x"0cff1151",
   132 => x"708025f2",
   133 => x"38bc0b86",
   134 => x"ffe19223",
   135 => x"81d40b86",
   136 => x"ffe19423",
   137 => x"80d9810b",
   138 => x"86ffe18e",
   139 => x"23e9c10b",
   140 => x"86ffe190",
   141 => x"2386ff0b",
   142 => x"86ffe380",
   143 => x"239fff0b",
   144 => x"86ffe382",
   145 => x"2381e00b",
   146 => x"8183a023",
   147 => x"81a00b90",
   148 => x"2c517081",
   149 => x"83a22381",
   150 => x"e20b8183",
   151 => x"a4237281",
   152 => x"83a623ff",
   153 => x"0b8183a8",
   154 => x"23fe0b81",
   155 => x"83aa2381",
   156 => x"83a00b90",
   157 => x"2c527186",
   158 => x"ffe18023",
   159 => x"8183a051",
   160 => x"7086ffe1",
   161 => x"8223800b",
   162 => x"86ffe188",
   163 => x"23fe8790",
   164 => x"0b86ffe1",
   165 => x"9623800b",
   166 => x"8183b00c",
   167 => x"800b8183",
   168 => x"b40c980b",
   169 => x"8183b80c",
   170 => x"028c050d",
   171 => x"0402f805",
   172 => x"0d8183b4",
   173 => x"08101081",
   174 => x"83b40805",
   175 => x"70902981",
   176 => x"83b00805",
   177 => x"85d01151",
   178 => x"52528052",
   179 => x"71713471",
   180 => x"81123471",
   181 => x"82123471",
   182 => x"83123480",
   183 => x"d0118113",
   184 => x"535181ff",
   185 => x"7225e538",
   186 => x"0288050d",
   187 => x"0402f405",
   188 => x"0d81a053",
   189 => x"a0bf5272",
   190 => x"84147108",
   191 => x"8105720c",
   192 => x"ff145454",
   193 => x"51807224",
   194 => x"e8387284",
   195 => x"14710881",
   196 => x"05720cff",
   197 => x"14545451",
   198 => x"718025db",
   199 => x"38a08085",
   200 => x"f10402e8",
   201 => x"050d7756",
   202 => x"9f762581",
   203 => x"90388183",
   204 => x"b4087010",
   205 => x"10117081",
   206 => x"80298183",
   207 => x"b0080585",
   208 => x"d0117910",
   209 => x"1010a080",
   210 => x"8a8c0570",
   211 => x"70840552",
   212 => x"08710852",
   213 => x"54555154",
   214 => x"55557072",
   215 => x"3470882c",
   216 => x"5372ffb0",
   217 => x"13347090",
   218 => x"2c5372fe",
   219 => x"e0133470",
   220 => x"982c5170",
   221 => x"fe901334",
   222 => x"73fdc013",
   223 => x"3473882c",
   224 => x"5372fcf0",
   225 => x"13347390",
   226 => x"2c5170fc",
   227 => x"a0133473",
   228 => x"982c5473",
   229 => x"fbd01334",
   230 => x"758a2eae",
   231 => x"388183b0",
   232 => x"08810581",
   233 => x"83b00c81",
   234 => x"83b00880",
   235 => x"d02e9b38",
   236 => x"74992eaf",
   237 => x"3875800c",
   238 => x"0298050d",
   239 => x"048183b4",
   240 => x"0855758a",
   241 => x"2e098106",
   242 => x"d4388115",
   243 => x"8183b40c",
   244 => x"800b8183",
   245 => x"b00c8183",
   246 => x"b4085574",
   247 => x"992e0981",
   248 => x"06d33881",
   249 => x"a00b8580",
   250 => x"118183b8",
   251 => x"08810581",
   252 => x"83b80c54",
   253 => x"528183b8",
   254 => x"08992ea6",
   255 => x"389f9f51",
   256 => x"72708405",
   257 => x"54087270",
   258 => x"8405540c",
   259 => x"ff115170",
   260 => x"8025ed38",
   261 => x"980b8183",
   262 => x"b40c7580",
   263 => x"0c029805",
   264 => x"0d0485ff",
   265 => x"c0813370",
   266 => x"862a8106",
   267 => x"515170f2",
   268 => x"38708183",
   269 => x"b80c9f9f",
   270 => x"51a08088",
   271 => x"800402d8",
   272 => x"050d7b59",
   273 => x"78708405",
   274 => x"5a085780",
   275 => x"5a76982a",
   276 => x"77882b58",
   277 => x"5675802e",
   278 => x"819e389f",
   279 => x"762581a0",
   280 => x"388183b4",
   281 => x"08701010",
   282 => x"11708180",
   283 => x"298183b0",
   284 => x"080585d0",
   285 => x"11791010",
   286 => x"10a0808a",
   287 => x"8c057070",
   288 => x"84055208",
   289 => x"71085254",
   290 => x"55515455",
   291 => x"55707234",
   292 => x"70882c53",
   293 => x"72ffb013",
   294 => x"3470902c",
   295 => x"5372fee0",
   296 => x"13347098",
   297 => x"2c5170fe",
   298 => x"90133473",
   299 => x"fdc01334",
   300 => x"73882c53",
   301 => x"72fcf013",
   302 => x"3473902c",
   303 => x"5170fca0",
   304 => x"13347398",
   305 => x"2c5473fb",
   306 => x"d0133475",
   307 => x"8a2ebe38",
   308 => x"8183b008",
   309 => x"81058183",
   310 => x"b00c8183",
   311 => x"b00880d0",
   312 => x"2eab3874",
   313 => x"992ebf38",
   314 => x"8118811b",
   315 => x"5b58837a",
   316 => x"25feda38",
   317 => x"75fecd38",
   318 => x"77800c02",
   319 => x"a8050d04",
   320 => x"8183b408",
   321 => x"55758a2e",
   322 => x"098106c4",
   323 => x"38811581",
   324 => x"83b40c80",
   325 => x"0b8183b0",
   326 => x"0c8183b4",
   327 => x"08557499",
   328 => x"2e098106",
   329 => x"c33881a0",
   330 => x"0b858011",
   331 => x"8183b808",
   332 => x"81058183",
   333 => x"b80c5452",
   334 => x"8183b808",
   335 => x"992eaf38",
   336 => x"9f9f5172",
   337 => x"70840554",
   338 => x"08727084",
   339 => x"05540cff",
   340 => x"11517080",
   341 => x"25ed3898",
   342 => x"0b8183b4",
   343 => x"0c811881",
   344 => x"1b5b5883",
   345 => x"7a25fde5",
   346 => x"38a08089",
   347 => x"f40485ff",
   348 => x"c0813370",
   349 => x"862a8106",
   350 => x"515170f2",
   351 => x"38708183",
   352 => x"b80c9f9f",
   353 => x"51a0808a",
   354 => x"c30402ec",
   355 => x"050d7654",
   356 => x"8755739c",
   357 => x"2a74842b",
   358 => x"b7125555",
   359 => x"52718924",
   360 => x"8438b012",
   361 => x"537251a0",
   362 => x"8086a22d",
   363 => x"ff155574",
   364 => x"8025df38",
   365 => x"0294050d",
   366 => x"0402f405",
   367 => x"0d830b85",
   368 => x"ffc48134",
   369 => x"fc0b85ff",
   370 => x"c08134a0",
   371 => x"8083d52d",
   372 => x"a0809a8c",
   373 => x"51a08088",
   374 => x"be2dff84",
   375 => x"0870892a",
   376 => x"70810651",
   377 => x"53537180",
   378 => x"2ef03872",
   379 => x"81ff0651",
   380 => x"a08086a2",
   381 => x"2da0808b",
   382 => x"da040000",
   383 => x"00ffffff",
   384 => x"ff00ffff",
   385 => x"ffff00ff",
   386 => x"ffffff00",
   387 => x"00000000",
   388 => x"00000000",
   389 => x"18181818",
   390 => x"18001800",
   391 => x"6c6c0000",
   392 => x"00000000",
   393 => x"6c6cfe6c",
   394 => x"fe6c6c00",
   395 => x"183e603c",
   396 => x"067c1800",
   397 => x"0066acd8",
   398 => x"366acc00",
   399 => x"386c6876",
   400 => x"dcce7b00",
   401 => x"18183000",
   402 => x"00000000",
   403 => x"0c183030",
   404 => x"30180c00",
   405 => x"30180c0c",
   406 => x"0c183000",
   407 => x"00663cff",
   408 => x"3c660000",
   409 => x"0018187e",
   410 => x"18180000",
   411 => x"00000000",
   412 => x"00181830",
   413 => x"0000007e",
   414 => x"00000000",
   415 => x"00000000",
   416 => x"00181800",
   417 => x"03060c18",
   418 => x"3060c000",
   419 => x"3c666e7e",
   420 => x"76663c00",
   421 => x"18387818",
   422 => x"18181800",
   423 => x"3c66060c",
   424 => x"18307e00",
   425 => x"3c66061c",
   426 => x"06663c00",
   427 => x"1c3c6ccc",
   428 => x"fe0c0c00",
   429 => x"7e607c06",
   430 => x"06663c00",
   431 => x"1c30607c",
   432 => x"66663c00",
   433 => x"7e06060c",
   434 => x"18181800",
   435 => x"3c66663c",
   436 => x"66663c00",
   437 => x"3c66663e",
   438 => x"060c3800",
   439 => x"00181800",
   440 => x"00181800",
   441 => x"00181800",
   442 => x"00181830",
   443 => x"00061860",
   444 => x"18060000",
   445 => x"00007e00",
   446 => x"7e000000",
   447 => x"00601806",
   448 => x"18600000",
   449 => x"3c66060c",
   450 => x"18001800",
   451 => x"7cc6ded6",
   452 => x"dec07800",
   453 => x"3c66667e",
   454 => x"66666600",
   455 => x"7c66667c",
   456 => x"66667c00",
   457 => x"1e306060",
   458 => x"60301e00",
   459 => x"786c6666",
   460 => x"666c7800",
   461 => x"7e606078",
   462 => x"60607e00",
   463 => x"7e606078",
   464 => x"60606000",
   465 => x"3c66606e",
   466 => x"66663e00",
   467 => x"6666667e",
   468 => x"66666600",
   469 => x"3c181818",
   470 => x"18183c00",
   471 => x"06060606",
   472 => x"06663c00",
   473 => x"c6ccd8f0",
   474 => x"d8ccc600",
   475 => x"60606060",
   476 => x"60607e00",
   477 => x"c6eefed6",
   478 => x"c6c6c600",
   479 => x"c6e6f6de",
   480 => x"cec6c600",
   481 => x"3c666666",
   482 => x"66663c00",
   483 => x"7c66667c",
   484 => x"60606000",
   485 => x"78cccccc",
   486 => x"ccdc7e00",
   487 => x"7c66667c",
   488 => x"6c666600",
   489 => x"3c66703c",
   490 => x"0e663c00",
   491 => x"7e181818",
   492 => x"18181800",
   493 => x"66666666",
   494 => x"66663c00",
   495 => x"66666666",
   496 => x"3c3c1800",
   497 => x"c6c6c6d6",
   498 => x"feeec600",
   499 => x"c3663c18",
   500 => x"3c66c300",
   501 => x"c3663c18",
   502 => x"18181800",
   503 => x"fe0c1830",
   504 => x"60c0fe00",
   505 => x"3c303030",
   506 => x"30303c00",
   507 => x"c0603018",
   508 => x"0c060300",
   509 => x"3c0c0c0c",
   510 => x"0c0c3c00",
   511 => x"10386cc6",
   512 => x"00000000",
   513 => x"00000000",
   514 => x"000000fe",
   515 => x"18180c00",
   516 => x"00000000",
   517 => x"00003c06",
   518 => x"3e663e00",
   519 => x"60607c66",
   520 => x"66667c00",
   521 => x"00003c60",
   522 => x"60603c00",
   523 => x"06063e66",
   524 => x"66663e00",
   525 => x"00003c66",
   526 => x"7e603c00",
   527 => x"1c307c30",
   528 => x"30303000",
   529 => x"00003e66",
   530 => x"663e063c",
   531 => x"60607c66",
   532 => x"66666600",
   533 => x"18001818",
   534 => x"18180c00",
   535 => x"0c000c0c",
   536 => x"0c0c0c78",
   537 => x"6060666c",
   538 => x"786c6600",
   539 => x"18181818",
   540 => x"18180c00",
   541 => x"0000ecfe",
   542 => x"d6c6c600",
   543 => x"00007c66",
   544 => x"66666600",
   545 => x"00003c66",
   546 => x"66663c00",
   547 => x"00007c66",
   548 => x"667c6060",
   549 => x"00003e66",
   550 => x"663e0606",
   551 => x"00007c66",
   552 => x"60606000",
   553 => x"00003c60",
   554 => x"3c067c00",
   555 => x"30307c30",
   556 => x"30301c00",
   557 => x"00006666",
   558 => x"66663e00",
   559 => x"00006666",
   560 => x"663c1800",
   561 => x"0000c6c6",
   562 => x"d6fe6c00",
   563 => x"0000c66c",
   564 => x"386cc600",
   565 => x"00006666",
   566 => x"663c1830",
   567 => x"00007e0c",
   568 => x"18307e00",
   569 => x"0e181870",
   570 => x"18180e00",
   571 => x"18181818",
   572 => x"18181800",
   573 => x"7018180e",
   574 => x"18187000",
   575 => x"729c0000",
   576 => x"00000000",
   577 => x"fefefefe",
   578 => x"fefefe00",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
   785 => x"00000000",
   786 => x"00000000",
   787 => x"00000000",
   788 => x"00000000",
   789 => x"00000000",
   790 => x"00000000",
   791 => x"00000000",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
   799 => x"00000000",
   800 => x"00000000",
   801 => x"00000000",
   802 => x"00000000",
   803 => x"00000000",
   804 => x"00000000",
   805 => x"00000000",
   806 => x"00000000",
   807 => x"00000000",
   808 => x"00000000",
   809 => x"00000000",
   810 => x"00000000",
   811 => x"00000000",
   812 => x"00000000",
   813 => x"00000000",
   814 => x"00000000",
   815 => x"00000000",
   816 => x"00000000",
   817 => x"00000000",
   818 => x"00000000",
   819 => x"00000000",
   820 => x"00000000",
   821 => x"00000000",
   822 => x"00000000",
   823 => x"00000000",
   824 => x"00000000",
   825 => x"00000000",
   826 => x"00000000",
   827 => x"00000000",
   828 => x"00000000",
   829 => x"00000000",
   830 => x"00000000",
   831 => x"00000000",
   832 => x"00000000",
   833 => x"00000000",
   834 => x"00000000",
   835 => x"52656164",
   836 => x"7920746f",
   837 => x"20726563",
   838 => x"65697665",
   839 => x"0a000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

