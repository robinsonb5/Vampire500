-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08081a3",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"89887383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02ec050d",
    30 => x"76548755",
    31 => x"739c2a74",
    32 => x"842bb712",
    33 => x"55555271",
    34 => x"89248438",
    35 => x"b0125372",
    36 => x"51a08084",
    37 => x"ae2dff15",
    38 => x"55748025",
    39 => x"df380294",
    40 => x"050d0402",
    41 => x"f4050d83",
    42 => x"0b85ffc4",
    43 => x"8134fc0b",
    44 => x"85ffc081",
    45 => x"34a08081",
    46 => x"e42da080",
    47 => x"899851a0",
    48 => x"8086c32d",
    49 => x"ff840870",
    50 => x"892a7081",
    51 => x"06515353",
    52 => x"71802ef0",
    53 => x"387281ff",
    54 => x"0651a080",
    55 => x"84ae2da0",
    56 => x"8081c404",
    57 => x"02f4050d",
    58 => x"fea0800b",
    59 => x"86ffe280",
    60 => x"23800b86",
    61 => x"ffe28223",
    62 => x"800b86ff",
    63 => x"e2842380",
    64 => x"0b86ffe2",
    65 => x"8823800b",
    66 => x"86ffe28a",
    67 => x"23907053",
    68 => x"53a0bf51",
    69 => x"80727084",
    70 => x"05540cff",
    71 => x"11517080",
    72 => x"25f238bc",
    73 => x"0b86ffe1",
    74 => x"922381d4",
    75 => x"0b86ffe1",
    76 => x"942380d9",
    77 => x"810b86ff",
    78 => x"e18e23e9",
    79 => x"c10b86ff",
    80 => x"e1902386",
    81 => x"ff0b86ff",
    82 => x"e380239f",
    83 => x"ff0b86ff",
    84 => x"e3822381",
    85 => x"e00b8182",
    86 => x"9023900b",
    87 => x"902c5170",
    88 => x"81829223",
    89 => x"81e20b81",
    90 => x"82942372",
    91 => x"81829623",
    92 => x"ff0b8182",
    93 => x"9823fe0b",
    94 => x"81829a23",
    95 => x"8182900b",
    96 => x"902c5271",
    97 => x"86ffe180",
    98 => x"23818290",
    99 => x"517086ff",
   100 => x"e1822380",
   101 => x"0b86ffe1",
   102 => x"8823fe87",
   103 => x"900b86ff",
   104 => x"e1962380",
   105 => x"0b8182a0",
   106 => x"0c800b81",
   107 => x"82a40c98",
   108 => x"0b8182a8",
   109 => x"0c028c05",
   110 => x"0d0402f8",
   111 => x"050d8182",
   112 => x"a4081010",
   113 => x"8182a408",
   114 => x"05709029",
   115 => x"8182a008",
   116 => x"0584c011",
   117 => x"51525280",
   118 => x"52717134",
   119 => x"71811234",
   120 => x"71821234",
   121 => x"71831234",
   122 => x"80d01181",
   123 => x"13535181",
   124 => x"ff7225e5",
   125 => x"38028805",
   126 => x"0d0402f4",
   127 => x"050d9053",
   128 => x"a0bf5272",
   129 => x"84147108",
   130 => x"8105720c",
   131 => x"ff145454",
   132 => x"51807224",
   133 => x"e9387284",
   134 => x"14710881",
   135 => x"05720cff",
   136 => x"14545451",
   137 => x"718025db",
   138 => x"38a08083",
   139 => x"fe0402e8",
   140 => x"050d7756",
   141 => x"9f762581",
   142 => x"8d388182",
   143 => x"a4087010",
   144 => x"10117081",
   145 => x"80298182",
   146 => x"a0080584",
   147 => x"c0117910",
   148 => x"1010a080",
   149 => x"87ac0570",
   150 => x"70840552",
   151 => x"08710852",
   152 => x"54555154",
   153 => x"55557072",
   154 => x"3470882c",
   155 => x"5372ffb0",
   156 => x"13347090",
   157 => x"2c5372fe",
   158 => x"e0133470",
   159 => x"982c5170",
   160 => x"fe901334",
   161 => x"73fdc013",
   162 => x"3473882c",
   163 => x"5372fcf0",
   164 => x"13347390",
   165 => x"2c5170fc",
   166 => x"a0133473",
   167 => x"982c5473",
   168 => x"fbd01334",
   169 => x"758a2eab",
   170 => x"388182a0",
   171 => x"08810581",
   172 => x"82a00c81",
   173 => x"82a00880",
   174 => x"d02e9838",
   175 => x"74992eac",
   176 => x"38029805",
   177 => x"0d048182",
   178 => x"a4085575",
   179 => x"8a2e0981",
   180 => x"06d73881",
   181 => x"158182a4",
   182 => x"0c800b81",
   183 => x"82a00c81",
   184 => x"82a40855",
   185 => x"74992e09",
   186 => x"8106d638",
   187 => x"900b8580",
   188 => x"118182a8",
   189 => x"08810581",
   190 => x"82a80c54",
   191 => x"528182a8",
   192 => x"08992ea3",
   193 => x"389f9f51",
   194 => x"72708405",
   195 => x"54087270",
   196 => x"8405540c",
   197 => x"ff115170",
   198 => x"8025ed38",
   199 => x"980b8182",
   200 => x"a40c0298",
   201 => x"050d0485",
   202 => x"ffc08133",
   203 => x"70862a81",
   204 => x"06525670",
   205 => x"f2387081",
   206 => x"82a80c9f",
   207 => x"9f51a080",
   208 => x"86880402",
   209 => x"dc050d7a",
   210 => x"58777084",
   211 => x"05590857",
   212 => x"80597698",
   213 => x"2a77882b",
   214 => x"58567580",
   215 => x"2e819b38",
   216 => x"9f762581",
   217 => x"9a388182",
   218 => x"a4087010",
   219 => x"10117081",
   220 => x"80298182",
   221 => x"a0080584",
   222 => x"c0117910",
   223 => x"1010a080",
   224 => x"87ac0570",
   225 => x"70840552",
   226 => x"08710852",
   227 => x"54555154",
   228 => x"55557072",
   229 => x"3470882c",
   230 => x"5372ffb0",
   231 => x"13347090",
   232 => x"2c5372fe",
   233 => x"e0133470",
   234 => x"982c5170",
   235 => x"fe901334",
   236 => x"73fdc013",
   237 => x"3473882c",
   238 => x"5372fcf0",
   239 => x"13347390",
   240 => x"2c5170fc",
   241 => x"a0133473",
   242 => x"982c5473",
   243 => x"fbd01334",
   244 => x"758a2eb8",
   245 => x"388182a0",
   246 => x"08810581",
   247 => x"82a00c81",
   248 => x"82a00880",
   249 => x"d02ea538",
   250 => x"74992eb9",
   251 => x"38811959",
   252 => x"837925fe",
   253 => x"dd3875fe",
   254 => x"d03802a4",
   255 => x"050d0481",
   256 => x"82a40855",
   257 => x"758a2e09",
   258 => x"8106ca38",
   259 => x"81158182",
   260 => x"a40c800b",
   261 => x"8182a00c",
   262 => x"8182a408",
   263 => x"5574992e",
   264 => x"098106c9",
   265 => x"38900b85",
   266 => x"80118182",
   267 => x"a8088105",
   268 => x"8182a80c",
   269 => x"54528182",
   270 => x"a808992e",
   271 => x"ac389f9f",
   272 => x"51727084",
   273 => x"05540872",
   274 => x"70840554",
   275 => x"0cff1151",
   276 => x"708025ed",
   277 => x"38980b81",
   278 => x"82a40c81",
   279 => x"19598379",
   280 => x"25fdef38",
   281 => x"a08087f6",
   282 => x"0485ffc0",
   283 => x"81337086",
   284 => x"2a810651",
   285 => x"5170f238",
   286 => x"708182a8",
   287 => x"0c9f9f51",
   288 => x"a08088c1",
   289 => x"04000000",
   290 => x"00ffffff",
   291 => x"ff00ffff",
   292 => x"ffff00ff",
   293 => x"ffffff00",
   294 => x"52656164",
   295 => x"7920746f",
   296 => x"20726563",
   297 => x"65697665",
   298 => x"0a000000",
   299 => x"00000000",
   300 => x"00000000",
   301 => x"18181818",
   302 => x"18001800",
   303 => x"6c6c0000",
   304 => x"00000000",
   305 => x"6c6cfe6c",
   306 => x"fe6c6c00",
   307 => x"183e603c",
   308 => x"067c1800",
   309 => x"0066acd8",
   310 => x"366acc00",
   311 => x"386c6876",
   312 => x"dcce7b00",
   313 => x"18183000",
   314 => x"00000000",
   315 => x"0c183030",
   316 => x"30180c00",
   317 => x"30180c0c",
   318 => x"0c183000",
   319 => x"00663cff",
   320 => x"3c660000",
   321 => x"0018187e",
   322 => x"18180000",
   323 => x"00000000",
   324 => x"00181830",
   325 => x"0000007e",
   326 => x"00000000",
   327 => x"00000000",
   328 => x"00181800",
   329 => x"03060c18",
   330 => x"3060c000",
   331 => x"3c666e7e",
   332 => x"76663c00",
   333 => x"18387818",
   334 => x"18181800",
   335 => x"3c66060c",
   336 => x"18307e00",
   337 => x"3c66061c",
   338 => x"06663c00",
   339 => x"1c3c6ccc",
   340 => x"fe0c0c00",
   341 => x"7e607c06",
   342 => x"06663c00",
   343 => x"1c30607c",
   344 => x"66663c00",
   345 => x"7e06060c",
   346 => x"18181800",
   347 => x"3c66663c",
   348 => x"66663c00",
   349 => x"3c66663e",
   350 => x"060c3800",
   351 => x"00181800",
   352 => x"00181800",
   353 => x"00181800",
   354 => x"00181830",
   355 => x"00061860",
   356 => x"18060000",
   357 => x"00007e00",
   358 => x"7e000000",
   359 => x"00601806",
   360 => x"18600000",
   361 => x"3c66060c",
   362 => x"18001800",
   363 => x"7cc6ded6",
   364 => x"dec07800",
   365 => x"3c66667e",
   366 => x"66666600",
   367 => x"7c66667c",
   368 => x"66667c00",
   369 => x"1e306060",
   370 => x"60301e00",
   371 => x"786c6666",
   372 => x"666c7800",
   373 => x"7e606078",
   374 => x"60607e00",
   375 => x"7e606078",
   376 => x"60606000",
   377 => x"3c66606e",
   378 => x"66663e00",
   379 => x"6666667e",
   380 => x"66666600",
   381 => x"3c181818",
   382 => x"18183c00",
   383 => x"06060606",
   384 => x"06663c00",
   385 => x"c6ccd8f0",
   386 => x"d8ccc600",
   387 => x"60606060",
   388 => x"60607e00",
   389 => x"c6eefed6",
   390 => x"c6c6c600",
   391 => x"c6e6f6de",
   392 => x"cec6c600",
   393 => x"3c666666",
   394 => x"66663c00",
   395 => x"7c66667c",
   396 => x"60606000",
   397 => x"78cccccc",
   398 => x"ccdc7e00",
   399 => x"7c66667c",
   400 => x"6c666600",
   401 => x"3c66703c",
   402 => x"0e663c00",
   403 => x"7e181818",
   404 => x"18181800",
   405 => x"66666666",
   406 => x"66663c00",
   407 => x"66666666",
   408 => x"3c3c1800",
   409 => x"c6c6c6d6",
   410 => x"feeec600",
   411 => x"c3663c18",
   412 => x"3c66c300",
   413 => x"c3663c18",
   414 => x"18181800",
   415 => x"fe0c1830",
   416 => x"60c0fe00",
   417 => x"3c303030",
   418 => x"30303c00",
   419 => x"c0603018",
   420 => x"0c060300",
   421 => x"3c0c0c0c",
   422 => x"0c0c3c00",
   423 => x"10386cc6",
   424 => x"00000000",
   425 => x"00000000",
   426 => x"000000fe",
   427 => x"18180c00",
   428 => x"00000000",
   429 => x"00003c06",
   430 => x"3e663e00",
   431 => x"60607c66",
   432 => x"66667c00",
   433 => x"00003c60",
   434 => x"60603c00",
   435 => x"06063e66",
   436 => x"66663e00",
   437 => x"00003c66",
   438 => x"7e603c00",
   439 => x"1c307c30",
   440 => x"30303000",
   441 => x"00003e66",
   442 => x"663e063c",
   443 => x"60607c66",
   444 => x"66666600",
   445 => x"18001818",
   446 => x"18180c00",
   447 => x"0c000c0c",
   448 => x"0c0c0c78",
   449 => x"6060666c",
   450 => x"786c6600",
   451 => x"18181818",
   452 => x"18180c00",
   453 => x"0000ecfe",
   454 => x"d6c6c600",
   455 => x"00007c66",
   456 => x"66666600",
   457 => x"00003c66",
   458 => x"66663c00",
   459 => x"00007c66",
   460 => x"667c6060",
   461 => x"00003e66",
   462 => x"663e0606",
   463 => x"00007c66",
   464 => x"60606000",
   465 => x"00003c60",
   466 => x"3c067c00",
   467 => x"30307c30",
   468 => x"30301c00",
   469 => x"00006666",
   470 => x"66663e00",
   471 => x"00006666",
   472 => x"663c1800",
   473 => x"0000c6c6",
   474 => x"d6fe6c00",
   475 => x"0000c66c",
   476 => x"386cc600",
   477 => x"00006666",
   478 => x"663c1830",
   479 => x"00007e0c",
   480 => x"18307e00",
   481 => x"0e181870",
   482 => x"18180e00",
   483 => x"18181818",
   484 => x"18181800",
   485 => x"7018180e",
   486 => x"18187000",
   487 => x"729c0000",
   488 => x"00000000",
   489 => x"fefefefe",
   490 => x"fefefe00",
   491 => x"00000000",
   492 => x"00000000",
   493 => x"00000000",
   494 => x"00000000",
   495 => x"00000000",
   496 => x"00000000",
   497 => x"00000000",
   498 => x"00000000",
   499 => x"00000000",
   500 => x"00000000",
   501 => x"00000000",
   502 => x"00000000",
   503 => x"00000000",
   504 => x"00000000",
   505 => x"00000000",
   506 => x"00000000",
   507 => x"00000000",
   508 => x"00000000",
   509 => x"00000000",
   510 => x"00000000",
   511 => x"00000000",
   512 => x"00000000",
   513 => x"00000000",
   514 => x"00000000",
   515 => x"00000000",
   516 => x"00000000",
   517 => x"00000000",
   518 => x"00000000",
   519 => x"00000000",
   520 => x"00000000",
   521 => x"00000000",
   522 => x"00000000",
   523 => x"00000000",
   524 => x"00000000",
   525 => x"00000000",
   526 => x"00000000",
   527 => x"00000000",
   528 => x"00000000",
   529 => x"00000000",
   530 => x"00000000",
   531 => x"00000000",
   532 => x"00000000",
   533 => x"00000000",
   534 => x"00000000",
   535 => x"00000000",
   536 => x"00000000",
   537 => x"00000000",
   538 => x"00000000",
   539 => x"00000000",
   540 => x"00000000",
   541 => x"00000000",
   542 => x"00000000",
   543 => x"00000000",
   544 => x"00000000",
   545 => x"00000000",
   546 => x"00000000",
   547 => x"00000000",
   548 => x"00000000",
   549 => x"00000000",
   550 => x"00000000",
   551 => x"00000000",
   552 => x"00000000",
   553 => x"00000000",
   554 => x"00000000",
   555 => x"00000000",
   556 => x"00000000",
   557 => x"00000000",
   558 => x"00000000",
   559 => x"00000000",
   560 => x"00000000",
   561 => x"00000000",
   562 => x"00000000",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

