-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08080f4",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"81987383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02f4050d",
    30 => x"80537281",
    31 => x"14545271",
    32 => x"86ffe380",
    33 => x"23728114",
    34 => x"54527186",
    35 => x"ffe38023",
    36 => x"a08080fa",
    37 => x"04000000",
    38 => x"00ffffff",
    39 => x"ff00ffff",
    40 => x"ffff00ff",
    41 => x"ffffff00",
    42 => x"00000000",
    43 => x"00000000",
    44 => x"18181818",
    45 => x"18001800",
    46 => x"6c6c0000",
    47 => x"00000000",
    48 => x"6c6cfe6c",
    49 => x"fe6c6c00",
    50 => x"183e603c",
    51 => x"067c1800",
    52 => x"0066acd8",
    53 => x"366acc00",
    54 => x"386c6876",
    55 => x"dcce7b00",
    56 => x"18183000",
    57 => x"00000000",
    58 => x"0c183030",
    59 => x"30180c00",
    60 => x"30180c0c",
    61 => x"0c183000",
    62 => x"00663cff",
    63 => x"3c660000",
    64 => x"0018187e",
    65 => x"18180000",
    66 => x"00000000",
    67 => x"00181830",
    68 => x"0000007e",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00181800",
    72 => x"03060c18",
    73 => x"3060c000",
    74 => x"3c666e7e",
    75 => x"76663c00",
    76 => x"18387818",
    77 => x"18181800",
    78 => x"3c66060c",
    79 => x"18307e00",
    80 => x"3c66061c",
    81 => x"06663c00",
    82 => x"1c3c6ccc",
    83 => x"fe0c0c00",
    84 => x"7e607c06",
    85 => x"06663c00",
    86 => x"1c30607c",
    87 => x"66663c00",
    88 => x"7e06060c",
    89 => x"18181800",
    90 => x"3c66663c",
    91 => x"66663c00",
    92 => x"3c66663e",
    93 => x"060c3800",
    94 => x"00181800",
    95 => x"00181800",
    96 => x"00181800",
    97 => x"00181830",
    98 => x"00061860",
    99 => x"18060000",
   100 => x"00007e00",
   101 => x"7e000000",
   102 => x"00601806",
   103 => x"18600000",
   104 => x"3c66060c",
   105 => x"18001800",
   106 => x"7cc6ded6",
   107 => x"dec07800",
   108 => x"3c66667e",
   109 => x"66666600",
   110 => x"7c66667c",
   111 => x"66667c00",
   112 => x"1e306060",
   113 => x"60301e00",
   114 => x"786c6666",
   115 => x"666c7800",
   116 => x"7e606078",
   117 => x"60607e00",
   118 => x"7e606078",
   119 => x"60606000",
   120 => x"3c66606e",
   121 => x"66663e00",
   122 => x"6666667e",
   123 => x"66666600",
   124 => x"3c181818",
   125 => x"18183c00",
   126 => x"06060606",
   127 => x"06663c00",
   128 => x"c6ccd8f0",
   129 => x"d8ccc600",
   130 => x"60606060",
   131 => x"60607e00",
   132 => x"c6eefed6",
   133 => x"c6c6c600",
   134 => x"c6e6f6de",
   135 => x"cec6c600",
   136 => x"3c666666",
   137 => x"66663c00",
   138 => x"7c66667c",
   139 => x"60606000",
   140 => x"78cccccc",
   141 => x"ccdc7e00",
   142 => x"7c66667c",
   143 => x"6c666600",
   144 => x"3c66703c",
   145 => x"0e663c00",
   146 => x"7e181818",
   147 => x"18181800",
   148 => x"66666666",
   149 => x"66663c00",
   150 => x"66666666",
   151 => x"3c3c1800",
   152 => x"c6c6c6d6",
   153 => x"feeec600",
   154 => x"c3663c18",
   155 => x"3c66c300",
   156 => x"c3663c18",
   157 => x"18181800",
   158 => x"fe0c1830",
   159 => x"60c0fe00",
   160 => x"3c303030",
   161 => x"30303c00",
   162 => x"c0603018",
   163 => x"0c060300",
   164 => x"3c0c0c0c",
   165 => x"0c0c3c00",
   166 => x"10386cc6",
   167 => x"00000000",
   168 => x"00000000",
   169 => x"000000fe",
   170 => x"18180c00",
   171 => x"00000000",
   172 => x"00003c06",
   173 => x"3e663e00",
   174 => x"60607c66",
   175 => x"66667c00",
   176 => x"00003c60",
   177 => x"60603c00",
   178 => x"06063e66",
   179 => x"66663e00",
   180 => x"00003c66",
   181 => x"7e603c00",
   182 => x"1c307c30",
   183 => x"30303000",
   184 => x"00003e66",
   185 => x"663e063c",
   186 => x"60607c66",
   187 => x"66666600",
   188 => x"18001818",
   189 => x"18180c00",
   190 => x"0c000c0c",
   191 => x"0c0c0c78",
   192 => x"6060666c",
   193 => x"786c6600",
   194 => x"18181818",
   195 => x"18180c00",
   196 => x"0000ecfe",
   197 => x"d6c6c600",
   198 => x"00007c66",
   199 => x"66666600",
   200 => x"00003c66",
   201 => x"66663c00",
   202 => x"00007c66",
   203 => x"667c6060",
   204 => x"00003e66",
   205 => x"663e0606",
   206 => x"00007c66",
   207 => x"60606000",
   208 => x"00003c60",
   209 => x"3c067c00",
   210 => x"30307c30",
   211 => x"30301c00",
   212 => x"00006666",
   213 => x"66663e00",
   214 => x"00006666",
   215 => x"663c1800",
   216 => x"0000c6c6",
   217 => x"d6fe6c00",
   218 => x"0000c66c",
   219 => x"386cc600",
   220 => x"00006666",
   221 => x"663c1830",
   222 => x"00007e0c",
   223 => x"18307e00",
   224 => x"0e181870",
   225 => x"18180e00",
   226 => x"18181818",
   227 => x"18181800",
   228 => x"7018180e",
   229 => x"18187000",
   230 => x"729c0000",
   231 => x"00000000",
   232 => x"fefefefe",
   233 => x"fefefe00",
   234 => x"00000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"00000000",
   249 => x"00000000",
   250 => x"00000000",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"00000000",
   257 => x"00000000",
   258 => x"00000000",
   259 => x"00000000",
   260 => x"00000000",
   261 => x"00000000",
   262 => x"00000000",
   263 => x"00000000",
   264 => x"00000000",
   265 => x"00000000",
   266 => x"00000000",
   267 => x"00000000",
   268 => x"00000000",
   269 => x"00000000",
   270 => x"00000000",
   271 => x"00000000",
   272 => x"00000000",
   273 => x"00000000",
   274 => x"00000000",
   275 => x"00000000",
   276 => x"00000000",
   277 => x"00000000",
   278 => x"00000000",
   279 => x"00000000",
   280 => x"00000000",
   281 => x"00000000",
   282 => x"00000000",
   283 => x"00000000",
   284 => x"00000000",
   285 => x"00000000",
   286 => x"00000000",
   287 => x"00000000",
   288 => x"00000000",
   289 => x"00000000",
   290 => x"00000000",
   291 => x"00000000",
   292 => x"00000000",
   293 => x"00000000",
   294 => x"00000000",
   295 => x"00000000",
   296 => x"00000000",
   297 => x"00000000",
   298 => x"00000000",
   299 => x"00000000",
   300 => x"00000000",
   301 => x"00000000",
   302 => x"00000000",
   303 => x"00000000",
   304 => x"00000000",
   305 => x"00000000",
   306 => x"00000000",
   307 => x"00000000",
   308 => x"00000000",
   309 => x"00000000",
   310 => x"00000000",
   311 => x"00000000",
   312 => x"00000000",
   313 => x"00000000",
   314 => x"00000000",
   315 => x"00000000",
   316 => x"00000000",
   317 => x"00000000",
   318 => x"00000000",
   319 => x"00000000",
   320 => x"00000000",
   321 => x"00000000",
   322 => x"00000000",
   323 => x"00000000",
   324 => x"00000000",
   325 => x"00000000",
   326 => x"00000000",
   327 => x"00000000",
   328 => x"00000000",
   329 => x"00000000",
   330 => x"00000000",
   331 => x"00000000",
   332 => x"00000000",
   333 => x"00000000",
   334 => x"00000000",
   335 => x"00000000",
   336 => x"00000000",
   337 => x"00000000",
   338 => x"00000000",
   339 => x"00000000",
   340 => x"00000000",
   341 => x"00000000",
   342 => x"00000000",
   343 => x"00000000",
   344 => x"00000000",
   345 => x"00000000",
   346 => x"00000000",
   347 => x"00000000",
   348 => x"00000000",
   349 => x"00000000",
   350 => x"00000000",
   351 => x"00000000",
   352 => x"00000000",
   353 => x"00000000",
   354 => x"00000000",
   355 => x"00000000",
   356 => x"00000000",
   357 => x"00000000",
   358 => x"00000000",
   359 => x"00000000",
   360 => x"00000000",
   361 => x"00000000",
   362 => x"00000000",
   363 => x"00000000",
   364 => x"00000000",
   365 => x"00000000",
   366 => x"00000000",
   367 => x"00000000",
   368 => x"00000000",
   369 => x"00000000",
   370 => x"00000000",
   371 => x"00000000",
   372 => x"00000000",
   373 => x"00000000",
   374 => x"00000000",
   375 => x"00000000",
   376 => x"00000000",
   377 => x"00000000",
   378 => x"00000000",
   379 => x"00000000",
   380 => x"00000000",
   381 => x"00000000",
   382 => x"00000000",
   383 => x"00000000",
   384 => x"00000000",
   385 => x"00000000",
   386 => x"00000000",
   387 => x"00000000",
   388 => x"00000000",
   389 => x"00000000",
   390 => x"00000000",
   391 => x"00000000",
   392 => x"00000000",
   393 => x"00000000",
   394 => x"00000000",
   395 => x"00000000",
   396 => x"00000000",
   397 => x"00000000",
   398 => x"00000000",
   399 => x"00000000",
   400 => x"00000000",
   401 => x"00000000",
   402 => x"00000000",
   403 => x"00000000",
   404 => x"00000000",
   405 => x"00000000",
   406 => x"00000000",
   407 => x"00000000",
   408 => x"00000000",
   409 => x"00000000",
   410 => x"00000000",
   411 => x"00000000",
   412 => x"00000000",
   413 => x"00000000",
   414 => x"00000000",
   415 => x"00000000",
   416 => x"00000000",
   417 => x"00000000",
   418 => x"00000000",
   419 => x"00000000",
   420 => x"00000000",
   421 => x"00000000",
   422 => x"00000000",
   423 => x"00000000",
   424 => x"00000000",
   425 => x"00000000",
   426 => x"00000000",
   427 => x"00000000",
   428 => x"00000000",
   429 => x"00000000",
   430 => x"00000000",
   431 => x"00000000",
   432 => x"00000000",
   433 => x"00000000",
   434 => x"00000000",
   435 => x"00000000",
   436 => x"00000000",
   437 => x"00000000",
   438 => x"00000000",
   439 => x"00000000",
   440 => x"00000000",
   441 => x"00000000",
   442 => x"00000000",
   443 => x"00000000",
   444 => x"00000000",
   445 => x"00000000",
   446 => x"00000000",
   447 => x"00000000",
   448 => x"00000000",
   449 => x"00000000",
   450 => x"00000000",
   451 => x"00000000",
   452 => x"00000000",
   453 => x"00000000",
   454 => x"00000000",
   455 => x"00000000",
   456 => x"00000000",
   457 => x"00000000",
   458 => x"00000000",
   459 => x"00000000",
   460 => x"00000000",
   461 => x"00000000",
   462 => x"00000000",
   463 => x"00000000",
   464 => x"00000000",
   465 => x"00000000",
   466 => x"00000000",
   467 => x"00000000",
   468 => x"00000000",
   469 => x"00000000",
   470 => x"00000000",
   471 => x"00000000",
   472 => x"00000000",
   473 => x"00000000",
   474 => x"00000000",
   475 => x"00000000",
   476 => x"00000000",
   477 => x"00000000",
   478 => x"00000000",
   479 => x"00000000",
   480 => x"00000000",
   481 => x"00000000",
   482 => x"00000000",
   483 => x"00000000",
   484 => x"00000000",
   485 => x"00000000",
   486 => x"00000000",
   487 => x"00000000",
   488 => x"00000000",
   489 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

