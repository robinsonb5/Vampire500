-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"f2040000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"8bec7383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040ba0",
    29 => x"8080fd0b",
    30 => x"a0808baa",
    31 => x"040ba080",
    32 => x"80fd0402",
    33 => x"c0050d02",
    34 => x"80c40580",
    35 => x"e05c5c80",
    36 => x"7c708405",
    37 => x"5e08715f",
    38 => x"5f587d70",
    39 => x"84055f08",
    40 => x"57805a76",
    41 => x"982a7788",
    42 => x"2b585574",
    43 => x"802e828d",
    44 => x"387c802e",
    45 => x"bf38805d",
    46 => x"7480e42e",
    47 => x"81af3874",
    48 => x"80e42680",
    49 => x"e8387480",
    50 => x"e32e80c1",
    51 => x"38a551a0",
    52 => x"8086932d",
    53 => x"7451a080",
    54 => x"86932d82",
    55 => x"1858811a",
    56 => x"5a837a25",
    57 => x"ffbd3874",
    58 => x"ffb0387e",
    59 => x"800c0280",
    60 => x"c0050d04",
    61 => x"74a52e09",
    62 => x"81069a38",
    63 => x"810b811b",
    64 => x"5b5d837a",
    65 => x"25ff9c38",
    66 => x"a08081e7",
    67 => x"047b841d",
    68 => x"7108575d",
    69 => x"547451a0",
    70 => x"8086932d",
    71 => x"8118811b",
    72 => x"5b58837a",
    73 => x"25fefc38",
    74 => x"a08081e7",
    75 => x"047480f3",
    76 => x"2e098106",
    77 => x"ff97387b",
    78 => x"841d7108",
    79 => x"70545d5d",
    80 => x"53a08088",
    81 => x"af2d800b",
    82 => x"ff115452",
    83 => x"807225ff",
    84 => x"8d387a70",
    85 => x"81055c33",
    86 => x"705255a0",
    87 => x"8086932d",
    88 => x"811873ff",
    89 => x"15555358",
    90 => x"a08082cc",
    91 => x"047b841d",
    92 => x"71087f5c",
    93 => x"555d5287",
    94 => x"56729c2a",
    95 => x"73842b54",
    96 => x"5271802e",
    97 => x"83388159",
    98 => x"b7125471",
    99 => x"89248438",
   100 => x"b0125478",
   101 => x"9438ff16",
   102 => x"56758025",
   103 => x"dc38800b",
   104 => x"ff115452",
   105 => x"a08082cc",
   106 => x"047351a0",
   107 => x"8086932d",
   108 => x"ff165675",
   109 => x"8025c238",
   110 => x"a080839e",
   111 => x"0477800c",
   112 => x"0280c005",
   113 => x"0d0402f4",
   114 => x"050dfea0",
   115 => x"800b86ff",
   116 => x"e2802380",
   117 => x"0b86ffe2",
   118 => x"8223800b",
   119 => x"86ffe284",
   120 => x"23800b86",
   121 => x"ffe28823",
   122 => x"800b86ff",
   123 => x"e28a2381",
   124 => x"a0705353",
   125 => x"a0bf5180",
   126 => x"72708405",
   127 => x"540cff11",
   128 => x"51708025",
   129 => x"f238bc0b",
   130 => x"86ffe192",
   131 => x"2381d40b",
   132 => x"86ffe194",
   133 => x"2380d981",
   134 => x"0b86ffe1",
   135 => x"8e23e9c1",
   136 => x"0b86ffe1",
   137 => x"902386ff",
   138 => x"0b86ffe3",
   139 => x"80239fff",
   140 => x"0b86ffe3",
   141 => x"822381e0",
   142 => x"0b8183a0",
   143 => x"2381a00b",
   144 => x"902c5170",
   145 => x"8183a223",
   146 => x"81e20b81",
   147 => x"83a42372",
   148 => x"8183a623",
   149 => x"ff0b8183",
   150 => x"a823fe0b",
   151 => x"8183aa23",
   152 => x"8183a00b",
   153 => x"902c5271",
   154 => x"86ffe180",
   155 => x"238183a0",
   156 => x"517086ff",
   157 => x"e1822380",
   158 => x"0b86ffe1",
   159 => x"8823fe87",
   160 => x"900b86ff",
   161 => x"e1962380",
   162 => x"0b8183b0",
   163 => x"0c800b81",
   164 => x"83b40c98",
   165 => x"0b8183b8",
   166 => x"0c028c05",
   167 => x"0d0402f8",
   168 => x"050d8183",
   169 => x"b4081010",
   170 => x"8183b408",
   171 => x"05709029",
   172 => x"8183b008",
   173 => x"0585d011",
   174 => x"51525280",
   175 => x"52717134",
   176 => x"71811234",
   177 => x"71821234",
   178 => x"71831234",
   179 => x"80d01181",
   180 => x"13535181",
   181 => x"ff7225e5",
   182 => x"38028805",
   183 => x"0d0402f4",
   184 => x"050d81a0",
   185 => x"53a0bf52",
   186 => x"72841471",
   187 => x"08810572",
   188 => x"0cff1454",
   189 => x"54518072",
   190 => x"24e83872",
   191 => x"84147108",
   192 => x"8105720c",
   193 => x"ff145454",
   194 => x"51718025",
   195 => x"db38a080",
   196 => x"85e20402",
   197 => x"e8050d77",
   198 => x"569f7625",
   199 => x"81903881",
   200 => x"83b40870",
   201 => x"10101170",
   202 => x"81802981",
   203 => x"83b00805",
   204 => x"85d01179",
   205 => x"101010a0",
   206 => x"8089fc05",
   207 => x"70708405",
   208 => x"52087108",
   209 => x"52545551",
   210 => x"54555570",
   211 => x"72347088",
   212 => x"2c5372ff",
   213 => x"b0133470",
   214 => x"902c5372",
   215 => x"fee01334",
   216 => x"70982c51",
   217 => x"70fe9013",
   218 => x"3473fdc0",
   219 => x"13347388",
   220 => x"2c5372fc",
   221 => x"f0133473",
   222 => x"902c5170",
   223 => x"fca01334",
   224 => x"73982c54",
   225 => x"73fbd013",
   226 => x"34758a2e",
   227 => x"ae388183",
   228 => x"b0088105",
   229 => x"8183b00c",
   230 => x"8183b008",
   231 => x"80d02e9b",
   232 => x"3874992e",
   233 => x"af387580",
   234 => x"0c029805",
   235 => x"0d048183",
   236 => x"b4085575",
   237 => x"8a2e0981",
   238 => x"06d43881",
   239 => x"158183b4",
   240 => x"0c800b81",
   241 => x"83b00c81",
   242 => x"83b40855",
   243 => x"74992e09",
   244 => x"8106d338",
   245 => x"81a00b85",
   246 => x"80118183",
   247 => x"b8088105",
   248 => x"8183b80c",
   249 => x"54528183",
   250 => x"b808992e",
   251 => x"a6389f9f",
   252 => x"51727084",
   253 => x"05540872",
   254 => x"70840554",
   255 => x"0cff1151",
   256 => x"708025ed",
   257 => x"38980b81",
   258 => x"83b40c75",
   259 => x"800c0298",
   260 => x"050d0485",
   261 => x"ffc08133",
   262 => x"70862a81",
   263 => x"06515170",
   264 => x"f2387081",
   265 => x"83b80c9f",
   266 => x"9f51a080",
   267 => x"87f10402",
   268 => x"d8050d7b",
   269 => x"59787084",
   270 => x"055a0857",
   271 => x"805a7698",
   272 => x"2a77882b",
   273 => x"58567580",
   274 => x"2e819e38",
   275 => x"9f762581",
   276 => x"a0388183",
   277 => x"b4087010",
   278 => x"10117081",
   279 => x"80298183",
   280 => x"b0080585",
   281 => x"d0117910",
   282 => x"1010a080",
   283 => x"89fc0570",
   284 => x"70840552",
   285 => x"08710852",
   286 => x"54555154",
   287 => x"55557072",
   288 => x"3470882c",
   289 => x"5372ffb0",
   290 => x"13347090",
   291 => x"2c5372fe",
   292 => x"e0133470",
   293 => x"982c5170",
   294 => x"fe901334",
   295 => x"73fdc013",
   296 => x"3473882c",
   297 => x"5372fcf0",
   298 => x"13347390",
   299 => x"2c5170fc",
   300 => x"a0133473",
   301 => x"982c5473",
   302 => x"fbd01334",
   303 => x"758a2ebe",
   304 => x"388183b0",
   305 => x"08810581",
   306 => x"83b00c81",
   307 => x"83b00880",
   308 => x"d02eab38",
   309 => x"74992ebf",
   310 => x"38811881",
   311 => x"1b5b5883",
   312 => x"7a25feda",
   313 => x"3875fecd",
   314 => x"3877800c",
   315 => x"02a8050d",
   316 => x"048183b4",
   317 => x"0855758a",
   318 => x"2e098106",
   319 => x"c4388115",
   320 => x"8183b40c",
   321 => x"800b8183",
   322 => x"b00c8183",
   323 => x"b4085574",
   324 => x"992e0981",
   325 => x"06c33881",
   326 => x"a00b8580",
   327 => x"118183b8",
   328 => x"08810581",
   329 => x"83b80c54",
   330 => x"528183b8",
   331 => x"08992eaf",
   332 => x"389f9f51",
   333 => x"72708405",
   334 => x"54087270",
   335 => x"8405540c",
   336 => x"ff115170",
   337 => x"8025ed38",
   338 => x"980b8183",
   339 => x"b40c8118",
   340 => x"811b5b58",
   341 => x"837a25fd",
   342 => x"e538a080",
   343 => x"89e50485",
   344 => x"ffc08133",
   345 => x"70862a81",
   346 => x"06515170",
   347 => x"f2387081",
   348 => x"83b80c9f",
   349 => x"9f51a080",
   350 => x"8ab40402",
   351 => x"ec050d76",
   352 => x"54875573",
   353 => x"9c2a7484",
   354 => x"2bb71255",
   355 => x"55527189",
   356 => x"248438b0",
   357 => x"12537251",
   358 => x"a0808693",
   359 => x"2dff1555",
   360 => x"748025df",
   361 => x"38029405",
   362 => x"0d0402f4",
   363 => x"050d830b",
   364 => x"85ffc481",
   365 => x"34fc0b85",
   366 => x"ffc08134",
   367 => x"a08083c6",
   368 => x"2da08099",
   369 => x"fc51a080",
   370 => x"88af2dff",
   371 => x"84087089",
   372 => x"2a708106",
   373 => x"51535371",
   374 => x"802ef038",
   375 => x"7281ff06",
   376 => x"51a08086",
   377 => x"932da080",
   378 => x"8bcb0400",
   379 => x"00ffffff",
   380 => x"ff00ffff",
   381 => x"ffff00ff",
   382 => x"ffffff00",
   383 => x"00000000",
   384 => x"00000000",
   385 => x"18181818",
   386 => x"18001800",
   387 => x"6c6c0000",
   388 => x"00000000",
   389 => x"6c6cfe6c",
   390 => x"fe6c6c00",
   391 => x"183e603c",
   392 => x"067c1800",
   393 => x"0066acd8",
   394 => x"366acc00",
   395 => x"386c6876",
   396 => x"dcce7b00",
   397 => x"18183000",
   398 => x"00000000",
   399 => x"0c183030",
   400 => x"30180c00",
   401 => x"30180c0c",
   402 => x"0c183000",
   403 => x"00663cff",
   404 => x"3c660000",
   405 => x"0018187e",
   406 => x"18180000",
   407 => x"00000000",
   408 => x"00181830",
   409 => x"0000007e",
   410 => x"00000000",
   411 => x"00000000",
   412 => x"00181800",
   413 => x"03060c18",
   414 => x"3060c000",
   415 => x"3c666e7e",
   416 => x"76663c00",
   417 => x"18387818",
   418 => x"18181800",
   419 => x"3c66060c",
   420 => x"18307e00",
   421 => x"3c66061c",
   422 => x"06663c00",
   423 => x"1c3c6ccc",
   424 => x"fe0c0c00",
   425 => x"7e607c06",
   426 => x"06663c00",
   427 => x"1c30607c",
   428 => x"66663c00",
   429 => x"7e06060c",
   430 => x"18181800",
   431 => x"3c66663c",
   432 => x"66663c00",
   433 => x"3c66663e",
   434 => x"060c3800",
   435 => x"00181800",
   436 => x"00181800",
   437 => x"00181800",
   438 => x"00181830",
   439 => x"00061860",
   440 => x"18060000",
   441 => x"00007e00",
   442 => x"7e000000",
   443 => x"00601806",
   444 => x"18600000",
   445 => x"3c66060c",
   446 => x"18001800",
   447 => x"7cc6ded6",
   448 => x"dec07800",
   449 => x"3c66667e",
   450 => x"66666600",
   451 => x"7c66667c",
   452 => x"66667c00",
   453 => x"1e306060",
   454 => x"60301e00",
   455 => x"786c6666",
   456 => x"666c7800",
   457 => x"7e606078",
   458 => x"60607e00",
   459 => x"7e606078",
   460 => x"60606000",
   461 => x"3c66606e",
   462 => x"66663e00",
   463 => x"6666667e",
   464 => x"66666600",
   465 => x"3c181818",
   466 => x"18183c00",
   467 => x"06060606",
   468 => x"06663c00",
   469 => x"c6ccd8f0",
   470 => x"d8ccc600",
   471 => x"60606060",
   472 => x"60607e00",
   473 => x"c6eefed6",
   474 => x"c6c6c600",
   475 => x"c6e6f6de",
   476 => x"cec6c600",
   477 => x"3c666666",
   478 => x"66663c00",
   479 => x"7c66667c",
   480 => x"60606000",
   481 => x"78cccccc",
   482 => x"ccdc7e00",
   483 => x"7c66667c",
   484 => x"6c666600",
   485 => x"3c66703c",
   486 => x"0e663c00",
   487 => x"7e181818",
   488 => x"18181800",
   489 => x"66666666",
   490 => x"66663c00",
   491 => x"66666666",
   492 => x"3c3c1800",
   493 => x"c6c6c6d6",
   494 => x"feeec600",
   495 => x"c3663c18",
   496 => x"3c66c300",
   497 => x"c3663c18",
   498 => x"18181800",
   499 => x"fe0c1830",
   500 => x"60c0fe00",
   501 => x"3c303030",
   502 => x"30303c00",
   503 => x"c0603018",
   504 => x"0c060300",
   505 => x"3c0c0c0c",
   506 => x"0c0c3c00",
   507 => x"10386cc6",
   508 => x"00000000",
   509 => x"00000000",
   510 => x"000000fe",
   511 => x"18180c00",
   512 => x"00000000",
   513 => x"00003c06",
   514 => x"3e663e00",
   515 => x"60607c66",
   516 => x"66667c00",
   517 => x"00003c60",
   518 => x"60603c00",
   519 => x"06063e66",
   520 => x"66663e00",
   521 => x"00003c66",
   522 => x"7e603c00",
   523 => x"1c307c30",
   524 => x"30303000",
   525 => x"00003e66",
   526 => x"663e063c",
   527 => x"60607c66",
   528 => x"66666600",
   529 => x"18001818",
   530 => x"18180c00",
   531 => x"0c000c0c",
   532 => x"0c0c0c78",
   533 => x"6060666c",
   534 => x"786c6600",
   535 => x"18181818",
   536 => x"18180c00",
   537 => x"0000ecfe",
   538 => x"d6c6c600",
   539 => x"00007c66",
   540 => x"66666600",
   541 => x"00003c66",
   542 => x"66663c00",
   543 => x"00007c66",
   544 => x"667c6060",
   545 => x"00003e66",
   546 => x"663e0606",
   547 => x"00007c66",
   548 => x"60606000",
   549 => x"00003c60",
   550 => x"3c067c00",
   551 => x"30307c30",
   552 => x"30301c00",
   553 => x"00006666",
   554 => x"66663e00",
   555 => x"00006666",
   556 => x"663c1800",
   557 => x"0000c6c6",
   558 => x"d6fe6c00",
   559 => x"0000c66c",
   560 => x"386cc600",
   561 => x"00006666",
   562 => x"663c1830",
   563 => x"00007e0c",
   564 => x"18307e00",
   565 => x"0e181870",
   566 => x"18180e00",
   567 => x"18181818",
   568 => x"18181800",
   569 => x"7018180e",
   570 => x"18187000",
   571 => x"729c0000",
   572 => x"00000000",
   573 => x"fefefefe",
   574 => x"fefefe00",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
   785 => x"00000000",
   786 => x"00000000",
   787 => x"00000000",
   788 => x"00000000",
   789 => x"00000000",
   790 => x"00000000",
   791 => x"00000000",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
   799 => x"00000000",
   800 => x"00000000",
   801 => x"00000000",
   802 => x"00000000",
   803 => x"00000000",
   804 => x"00000000",
   805 => x"00000000",
   806 => x"00000000",
   807 => x"00000000",
   808 => x"00000000",
   809 => x"00000000",
   810 => x"00000000",
   811 => x"00000000",
   812 => x"00000000",
   813 => x"00000000",
   814 => x"00000000",
   815 => x"00000000",
   816 => x"00000000",
   817 => x"00000000",
   818 => x"00000000",
   819 => x"00000000",
   820 => x"00000000",
   821 => x"00000000",
   822 => x"00000000",
   823 => x"00000000",
   824 => x"00000000",
   825 => x"00000000",
   826 => x"00000000",
   827 => x"00000000",
   828 => x"00000000",
   829 => x"00000000",
   830 => x"00000000",
   831 => x"52656164",
   832 => x"7920746f",
   833 => x"20726563",
   834 => x"65697665",
   835 => x"0a000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

