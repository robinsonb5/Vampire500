SysClock_inst : SysClock PORT MAP (
		inclk0	 => inclk0_sig,
		pllena	 => pllena_sig,
		c0	 => c0_sig,
		c1	 => c1_sig
	);
