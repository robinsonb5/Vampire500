-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08080f4",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"87947383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02fc050d",
    30 => x"830b85ff",
    31 => x"c48134fc",
    32 => x"0b85ffc0",
    33 => x"8134a080",
    34 => x"81c92d80",
    35 => x"c851a080",
    36 => x"83992d80",
    37 => x"e551a080",
    38 => x"83992d80",
    39 => x"ec51a080",
    40 => x"83992d80",
    41 => x"ec51a080",
    42 => x"83992d80",
    43 => x"ef51a080",
    44 => x"83992d8a",
    45 => x"51a08083",
    46 => x"992da080",
    47 => x"87a451a0",
    48 => x"8084fe2d",
    49 => x"a08081c4",
    50 => x"0402f405",
    51 => x"0dfea080",
    52 => x"0b86ffe2",
    53 => x"8023800b",
    54 => x"86ffe282",
    55 => x"23800b86",
    56 => x"ffe28423",
    57 => x"800b86ff",
    58 => x"e2882380",
    59 => x"0b86ffe2",
    60 => x"8a239070",
    61 => x"5353a0bf",
    62 => x"51807270",
    63 => x"8405540c",
    64 => x"ff115170",
    65 => x"8025f238",
    66 => x"bc0b86ff",
    67 => x"e1922381",
    68 => x"d40b86ff",
    69 => x"e1942380",
    70 => x"d9810b86",
    71 => x"ffe18e23",
    72 => x"e9c10b86",
    73 => x"ffe19023",
    74 => x"86ff0b86",
    75 => x"ffe38023",
    76 => x"9fff0b86",
    77 => x"ffe38223",
    78 => x"81e00b84",
    79 => x"88902390",
    80 => x"0b902c51",
    81 => x"70848892",
    82 => x"2381e20b",
    83 => x"84889423",
    84 => x"72848896",
    85 => x"23ff0b84",
    86 => x"889823fe",
    87 => x"0b84889a",
    88 => x"23848890",
    89 => x"0b902c52",
    90 => x"7186ffe1",
    91 => x"80238488",
    92 => x"90517086",
    93 => x"ffe18223",
    94 => x"800b86ff",
    95 => x"e18823fe",
    96 => x"87900b86",
    97 => x"ffe19623",
    98 => x"800b8488",
    99 => x"a00c800b",
   100 => x"8488a40c",
   101 => x"028c050d",
   102 => x"0402e405",
   103 => x"0d02a305",
   104 => x"338488a4",
   105 => x"08701010",
   106 => x"118488a0",
   107 => x"08719029",
   108 => x"1184c011",
   109 => x"75a02917",
   110 => x"f8801108",
   111 => x"f8841208",
   112 => x"565a5751",
   113 => x"565a5657",
   114 => x"55727234",
   115 => x"72882c51",
   116 => x"70ffb013",
   117 => x"3472902c",
   118 => x"5170fee0",
   119 => x"13347298",
   120 => x"2c5170fe",
   121 => x"90133473",
   122 => x"fdc01334",
   123 => x"73882c53",
   124 => x"72fcf013",
   125 => x"3473902c",
   126 => x"5170fca0",
   127 => x"13347398",
   128 => x"2c5473fb",
   129 => x"d0133474",
   130 => x"8a2e80e2",
   131 => x"38811784",
   132 => x"88a00c84",
   133 => x"88a00880",
   134 => x"d02eb438",
   135 => x"75992e86",
   136 => x"38029c05",
   137 => x"0d04900b",
   138 => x"94801154",
   139 => x"529f9f51",
   140 => x"72708405",
   141 => x"54087270",
   142 => x"8405540c",
   143 => x"ff115170",
   144 => x"8025ed38",
   145 => x"980b8488",
   146 => x"a40c029c",
   147 => x"050d0481",
   148 => x"168488a4",
   149 => x"0c800b84",
   150 => x"88a00c84",
   151 => x"88a40856",
   152 => x"75992e09",
   153 => x"8106ffb9",
   154 => x"38a08084",
   155 => x"a6048116",
   156 => x"8488a40c",
   157 => x"8488a408",
   158 => x"56a08084",
   159 => x"e00402d4",
   160 => x"050d7c59",
   161 => x"78708405",
   162 => x"5a085780",
   163 => x"5a76982a",
   164 => x"77882b58",
   165 => x"5675802e",
   166 => x"81923884",
   167 => x"88a40870",
   168 => x"10101184",
   169 => x"88a00871",
   170 => x"90291184",
   171 => x"c0117aa0",
   172 => x"296005f8",
   173 => x"801108f8",
   174 => x"84120856",
   175 => x"59f88805",
   176 => x"4051555a",
   177 => x"55557272",
   178 => x"3472882c",
   179 => x"5170ffb0",
   180 => x"13347290",
   181 => x"2c5170fe",
   182 => x"e0133472",
   183 => x"982c5170",
   184 => x"fe901334",
   185 => x"73fdc013",
   186 => x"3473882c",
   187 => x"5372fcf0",
   188 => x"13347390",
   189 => x"2c5170fc",
   190 => x"a0133473",
   191 => x"982c5473",
   192 => x"fbd01334",
   193 => x"758a2e80",
   194 => x"f9388118",
   195 => x"8488a00c",
   196 => x"8488a008",
   197 => x"80d02e80",
   198 => x"ca387499",
   199 => x"2e933881",
   200 => x"1a5a837a",
   201 => x"25fee638",
   202 => x"75fed938",
   203 => x"02ac050d",
   204 => x"04900b94",
   205 => x"80115452",
   206 => x"9f9f5172",
   207 => x"70840554",
   208 => x"08727084",
   209 => x"05540cff",
   210 => x"11517080",
   211 => x"25ed3898",
   212 => x"0b8488a4",
   213 => x"0c811a5a",
   214 => x"837a25fe",
   215 => x"b038a080",
   216 => x"86a80481",
   217 => x"158488a4",
   218 => x"0c800b84",
   219 => x"88a00c84",
   220 => x"88a40855",
   221 => x"74992e09",
   222 => x"8106ffa3",
   223 => x"38a08086",
   224 => x"b1048115",
   225 => x"8488a40c",
   226 => x"8488a408",
   227 => x"55a08086",
   228 => x"f4040000",
   229 => x"00ffffff",
   230 => x"ff00ffff",
   231 => x"ffff00ff",
   232 => x"ffffff00",
   233 => x"48656c6c",
   234 => x"6f2c2077",
   235 => x"6f726c64",
   236 => x"210a0000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"18181818",
   240 => x"18001800",
   241 => x"6c6c0000",
   242 => x"00000000",
   243 => x"6c6cfe6c",
   244 => x"fe6c6c00",
   245 => x"183e603c",
   246 => x"067c1800",
   247 => x"0066acd8",
   248 => x"366acc00",
   249 => x"386c6876",
   250 => x"dcce7b00",
   251 => x"18183000",
   252 => x"00000000",
   253 => x"0c183030",
   254 => x"30180c00",
   255 => x"30180c0c",
   256 => x"0c183000",
   257 => x"00663cff",
   258 => x"3c660000",
   259 => x"0018187e",
   260 => x"18180000",
   261 => x"00000000",
   262 => x"00181830",
   263 => x"0000007e",
   264 => x"00000000",
   265 => x"00000000",
   266 => x"00181800",
   267 => x"03060c18",
   268 => x"3060c000",
   269 => x"3c666e7e",
   270 => x"76663c00",
   271 => x"18387818",
   272 => x"18181800",
   273 => x"3c66060c",
   274 => x"18307e00",
   275 => x"3c66061c",
   276 => x"06663c00",
   277 => x"1c3c6ccc",
   278 => x"fe0c0c00",
   279 => x"7e607c06",
   280 => x"06663c00",
   281 => x"1c30607c",
   282 => x"66663c00",
   283 => x"7e06060c",
   284 => x"18181800",
   285 => x"3c66663c",
   286 => x"66663c00",
   287 => x"3c66663e",
   288 => x"060c3800",
   289 => x"00181800",
   290 => x"00181800",
   291 => x"00181800",
   292 => x"00181830",
   293 => x"00061860",
   294 => x"18060000",
   295 => x"00007e00",
   296 => x"7e000000",
   297 => x"00601806",
   298 => x"18600000",
   299 => x"3c66060c",
   300 => x"18001800",
   301 => x"7cc6ded6",
   302 => x"dec07800",
   303 => x"3c66667e",
   304 => x"66666600",
   305 => x"7c66667c",
   306 => x"66667c00",
   307 => x"1e306060",
   308 => x"60301e00",
   309 => x"786c6666",
   310 => x"666c7800",
   311 => x"7e606078",
   312 => x"60607e00",
   313 => x"7e606078",
   314 => x"60606000",
   315 => x"3c66606e",
   316 => x"66663e00",
   317 => x"6666667e",
   318 => x"66666600",
   319 => x"3c181818",
   320 => x"18183c00",
   321 => x"06060606",
   322 => x"06663c00",
   323 => x"c6ccd8f0",
   324 => x"d8ccc600",
   325 => x"60606060",
   326 => x"60607e00",
   327 => x"c6eefed6",
   328 => x"c6c6c600",
   329 => x"c6e6f6de",
   330 => x"cec6c600",
   331 => x"3c666666",
   332 => x"66663c00",
   333 => x"7c66667c",
   334 => x"60606000",
   335 => x"78cccccc",
   336 => x"ccdc7e00",
   337 => x"7c66667c",
   338 => x"6c666600",
   339 => x"3c66703c",
   340 => x"0e663c00",
   341 => x"7e181818",
   342 => x"18181800",
   343 => x"66666666",
   344 => x"66663c00",
   345 => x"66666666",
   346 => x"3c3c1800",
   347 => x"c6c6c6d6",
   348 => x"feeec600",
   349 => x"c3663c18",
   350 => x"3c66c300",
   351 => x"c3663c18",
   352 => x"18181800",
   353 => x"fe0c1830",
   354 => x"60c0fe00",
   355 => x"3c303030",
   356 => x"30303c00",
   357 => x"c0603018",
   358 => x"0c060300",
   359 => x"3c0c0c0c",
   360 => x"0c0c3c00",
   361 => x"10386cc6",
   362 => x"00000000",
   363 => x"00000000",
   364 => x"000000fe",
   365 => x"18180c00",
   366 => x"00000000",
   367 => x"00003c06",
   368 => x"3e663e00",
   369 => x"60607c66",
   370 => x"66667c00",
   371 => x"00003c60",
   372 => x"60603c00",
   373 => x"06063e66",
   374 => x"66663e00",
   375 => x"00003c66",
   376 => x"7e603c00",
   377 => x"1c307c30",
   378 => x"30303000",
   379 => x"00003e66",
   380 => x"663e063c",
   381 => x"60607c66",
   382 => x"66666600",
   383 => x"18001818",
   384 => x"18180c00",
   385 => x"0c000c0c",
   386 => x"0c0c0c78",
   387 => x"6060666c",
   388 => x"786c6600",
   389 => x"18181818",
   390 => x"18180c00",
   391 => x"0000ecfe",
   392 => x"d6c6c600",
   393 => x"00007c66",
   394 => x"66666600",
   395 => x"00003c66",
   396 => x"66663c00",
   397 => x"00007c66",
   398 => x"667c6060",
   399 => x"00003e66",
   400 => x"663e0606",
   401 => x"00007c66",
   402 => x"60606000",
   403 => x"00003c60",
   404 => x"3c067c00",
   405 => x"30307c30",
   406 => x"30301c00",
   407 => x"00006666",
   408 => x"66663e00",
   409 => x"00006666",
   410 => x"663c1800",
   411 => x"0000c6c6",
   412 => x"d6fe6c00",
   413 => x"0000c66c",
   414 => x"386cc600",
   415 => x"00006666",
   416 => x"663c1830",
   417 => x"00007e0c",
   418 => x"18307e00",
   419 => x"0e181870",
   420 => x"18180e00",
   421 => x"18181818",
   422 => x"18181800",
   423 => x"7018180e",
   424 => x"18187000",
   425 => x"729c0000",
   426 => x"00000000",
   427 => x"fefefefe",
   428 => x"fefefe00",
   429 => x"00000000",
   430 => x"00000000",
   431 => x"00000000",
   432 => x"00000000",
   433 => x"00000000",
   434 => x"00000000",
   435 => x"00000000",
   436 => x"00000000",
   437 => x"00000000",
   438 => x"00000000",
   439 => x"00000000",
   440 => x"00000000",
   441 => x"00000000",
   442 => x"00000000",
   443 => x"00000000",
   444 => x"00000000",
   445 => x"00000000",
   446 => x"00000000",
   447 => x"00000000",
   448 => x"00000000",
   449 => x"00000000",
   450 => x"00000000",
   451 => x"00000000",
   452 => x"00000000",
   453 => x"00000000",
   454 => x"00000000",
   455 => x"00000000",
   456 => x"00000000",
   457 => x"00000000",
   458 => x"00000000",
   459 => x"00000000",
   460 => x"00000000",
   461 => x"00000000",
   462 => x"00000000",
   463 => x"00000000",
   464 => x"00000000",
   465 => x"00000000",
   466 => x"00000000",
   467 => x"00000000",
   468 => x"00000000",
   469 => x"00000000",
   470 => x"00000000",
   471 => x"00000000",
   472 => x"00000000",
   473 => x"00000000",
   474 => x"00000000",
   475 => x"00000000",
   476 => x"00000000",
   477 => x"00000000",
   478 => x"00000000",
   479 => x"00000000",
   480 => x"00000000",
   481 => x"00000000",
   482 => x"00000000",
   483 => x"00000000",
   484 => x"00000000",
   485 => x"00000000",
   486 => x"00000000",
   487 => x"00000000",
   488 => x"00000000",
   489 => x"00000000",
   490 => x"00000000",
   491 => x"00000000",
   492 => x"00000000",
   493 => x"00000000",
   494 => x"00000000",
   495 => x"00000000",
   496 => x"00000000",
   497 => x"00000000",
   498 => x"00000000",
   499 => x"00000000",
   500 => x"00000000",
   501 => x"00000000",
   502 => x"00000000",
   503 => x"00000000",
   504 => x"00000000",
   505 => x"00000000",
   506 => x"00000000",
   507 => x"00000000",
   508 => x"00000000",
   509 => x"00000000",
   510 => x"00000000",
   511 => x"00000000",
   512 => x"00000000",
   513 => x"00000000",
   514 => x"00000000",
   515 => x"00000000",
   516 => x"00000000",
   517 => x"00000000",
   518 => x"00000000",
   519 => x"00000000",
   520 => x"00000000",
   521 => x"00000000",
   522 => x"00000000",
   523 => x"00000000",
   524 => x"00000000",
   525 => x"00000000",
   526 => x"00000000",
   527 => x"00000000",
   528 => x"00000000",
   529 => x"00000000",
   530 => x"00000000",
   531 => x"00000000",
   532 => x"00000000",
   533 => x"00000000",
   534 => x"00000000",
   535 => x"00000000",
   536 => x"00000000",
   537 => x"00000000",
   538 => x"00000000",
   539 => x"00000000",
   540 => x"00000000",
   541 => x"00000000",
   542 => x"00000000",
   543 => x"00000000",
   544 => x"00000000",
   545 => x"00000000",
   546 => x"00000000",
   547 => x"00000000",
   548 => x"00000000",
   549 => x"00000000",
   550 => x"00000000",
   551 => x"00000000",
   552 => x"00000000",
   553 => x"00000000",
   554 => x"00000000",
   555 => x"00000000",
   556 => x"00000000",
   557 => x"00000000",
   558 => x"00000000",
   559 => x"00000000",
   560 => x"00000000",
   561 => x"00000000",
   562 => x"00000000",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

