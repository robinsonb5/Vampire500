-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08081a3",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"88a47383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02ec050d",
    30 => x"76548755",
    31 => x"739c2a74",
    32 => x"842bb712",
    33 => x"55555271",
    34 => x"89248438",
    35 => x"b0125372",
    36 => x"51a08084",
    37 => x"a82dff15",
    38 => x"55748025",
    39 => x"df380294",
    40 => x"050d0402",
    41 => x"f4050d83",
    42 => x"0b85ffc4",
    43 => x"8134fc0b",
    44 => x"85ffc081",
    45 => x"34a08081",
    46 => x"e42da080",
    47 => x"88b451a0",
    48 => x"80868f2d",
    49 => x"ff840870",
    50 => x"892a7081",
    51 => x"06515353",
    52 => x"71802ef0",
    53 => x"387281ff",
    54 => x"0651a080",
    55 => x"84a82da0",
    56 => x"8081c404",
    57 => x"02f4050d",
    58 => x"fea0800b",
    59 => x"86ffe280",
    60 => x"23800b86",
    61 => x"ffe28223",
    62 => x"800b86ff",
    63 => x"e2842380",
    64 => x"0b86ffe2",
    65 => x"8823800b",
    66 => x"86ffe28a",
    67 => x"23907053",
    68 => x"53a0bf51",
    69 => x"80727084",
    70 => x"05540cff",
    71 => x"11517080",
    72 => x"25f238bc",
    73 => x"0b86ffe1",
    74 => x"922381d4",
    75 => x"0b86ffe1",
    76 => x"942380d9",
    77 => x"810b86ff",
    78 => x"e18e23e9",
    79 => x"c10b86ff",
    80 => x"e1902386",
    81 => x"ff0b86ff",
    82 => x"e380239f",
    83 => x"ff0b86ff",
    84 => x"e3822381",
    85 => x"e00b8182",
    86 => x"9023900b",
    87 => x"902c5170",
    88 => x"81829223",
    89 => x"81e20b81",
    90 => x"82942372",
    91 => x"81829623",
    92 => x"ff0b8182",
    93 => x"9823fe0b",
    94 => x"81829a23",
    95 => x"8182900b",
    96 => x"902c5271",
    97 => x"86ffe180",
    98 => x"23818290",
    99 => x"517086ff",
   100 => x"e1822380",
   101 => x"0b86ffe1",
   102 => x"8823fe87",
   103 => x"900b86ff",
   104 => x"e1962380",
   105 => x"0b8182a0",
   106 => x"0c800b81",
   107 => x"82a40c02",
   108 => x"8c050d04",
   109 => x"02f8050d",
   110 => x"8182a408",
   111 => x"10108182",
   112 => x"a4080570",
   113 => x"90298182",
   114 => x"a0080584",
   115 => x"c0115152",
   116 => x"52805271",
   117 => x"71347181",
   118 => x"12347182",
   119 => x"12347183",
   120 => x"123480d0",
   121 => x"11811353",
   122 => x"5181ff72",
   123 => x"25e53802",
   124 => x"88050d04",
   125 => x"02f4050d",
   126 => x"9053a0bf",
   127 => x"52728414",
   128 => x"71088105",
   129 => x"720cff14",
   130 => x"54545180",
   131 => x"7224e938",
   132 => x"72841471",
   133 => x"08810572",
   134 => x"0cff1454",
   135 => x"54517180",
   136 => x"25db38a0",
   137 => x"8083f804",
   138 => x"02e8050d",
   139 => x"77569f76",
   140 => x"25818d38",
   141 => x"8182a408",
   142 => x"70101011",
   143 => x"70818029",
   144 => x"8182a008",
   145 => x"0584c011",
   146 => x"79101010",
   147 => x"a08086c8",
   148 => x"05707084",
   149 => x"05520871",
   150 => x"08525455",
   151 => x"51545555",
   152 => x"70723470",
   153 => x"882c5372",
   154 => x"ffb01334",
   155 => x"70902c53",
   156 => x"72fee013",
   157 => x"3470982c",
   158 => x"5170fe90",
   159 => x"133473fd",
   160 => x"c0133473",
   161 => x"882c5372",
   162 => x"fcf01334",
   163 => x"73902c51",
   164 => x"70fca013",
   165 => x"3473982c",
   166 => x"5473fbd0",
   167 => x"1334758a",
   168 => x"2eab3881",
   169 => x"82a00881",
   170 => x"058182a0",
   171 => x"0c8182a0",
   172 => x"0880d02e",
   173 => x"98387499",
   174 => x"2eac3802",
   175 => x"98050d04",
   176 => x"8182a408",
   177 => x"55758a2e",
   178 => x"098106d7",
   179 => x"38811581",
   180 => x"82a40c80",
   181 => x"0b8182a0",
   182 => x"0c8182a4",
   183 => x"08557499",
   184 => x"2e098106",
   185 => x"d638900b",
   186 => x"85801154",
   187 => x"529f9f51",
   188 => x"72708405",
   189 => x"54087270",
   190 => x"8405540c",
   191 => x"ff115170",
   192 => x"8025ed38",
   193 => x"980b8182",
   194 => x"a40c0298",
   195 => x"050d0402",
   196 => x"dc050d7a",
   197 => x"58777084",
   198 => x"05590857",
   199 => x"80597698",
   200 => x"2a77882b",
   201 => x"58567580",
   202 => x"2e819b38",
   203 => x"9f762581",
   204 => x"9a388182",
   205 => x"a4087010",
   206 => x"10117081",
   207 => x"80298182",
   208 => x"a0080584",
   209 => x"c0117910",
   210 => x"1010a080",
   211 => x"86c80570",
   212 => x"70840552",
   213 => x"08710852",
   214 => x"54555154",
   215 => x"55557072",
   216 => x"3470882c",
   217 => x"5372ffb0",
   218 => x"13347090",
   219 => x"2c5372fe",
   220 => x"e0133470",
   221 => x"982c5170",
   222 => x"fe901334",
   223 => x"73fdc013",
   224 => x"3473882c",
   225 => x"5372fcf0",
   226 => x"13347390",
   227 => x"2c5170fc",
   228 => x"a0133473",
   229 => x"982c5473",
   230 => x"fbd01334",
   231 => x"758a2eb8",
   232 => x"388182a0",
   233 => x"08810581",
   234 => x"82a00c81",
   235 => x"82a00880",
   236 => x"d02ea538",
   237 => x"74992eb9",
   238 => x"38811959",
   239 => x"837925fe",
   240 => x"dd3875fe",
   241 => x"d03802a4",
   242 => x"050d0481",
   243 => x"82a40855",
   244 => x"758a2e09",
   245 => x"8106ca38",
   246 => x"81158182",
   247 => x"a40c800b",
   248 => x"8182a00c",
   249 => x"8182a408",
   250 => x"5574992e",
   251 => x"098106c9",
   252 => x"38900b85",
   253 => x"80115452",
   254 => x"9f9f5172",
   255 => x"70840554",
   256 => x"08727084",
   257 => x"05540cff",
   258 => x"11517080",
   259 => x"25ed3898",
   260 => x"0b8182a4",
   261 => x"0c811959",
   262 => x"837925fe",
   263 => x"8138a080",
   264 => x"87c20400",
   265 => x"00ffffff",
   266 => x"ff00ffff",
   267 => x"ffff00ff",
   268 => x"ffffff00",
   269 => x"52656164",
   270 => x"7920746f",
   271 => x"20726563",
   272 => x"65697665",
   273 => x"0a000000",
   274 => x"00000000",
   275 => x"00000000",
   276 => x"18181818",
   277 => x"18001800",
   278 => x"6c6c0000",
   279 => x"00000000",
   280 => x"6c6cfe6c",
   281 => x"fe6c6c00",
   282 => x"183e603c",
   283 => x"067c1800",
   284 => x"0066acd8",
   285 => x"366acc00",
   286 => x"386c6876",
   287 => x"dcce7b00",
   288 => x"18183000",
   289 => x"00000000",
   290 => x"0c183030",
   291 => x"30180c00",
   292 => x"30180c0c",
   293 => x"0c183000",
   294 => x"00663cff",
   295 => x"3c660000",
   296 => x"0018187e",
   297 => x"18180000",
   298 => x"00000000",
   299 => x"00181830",
   300 => x"0000007e",
   301 => x"00000000",
   302 => x"00000000",
   303 => x"00181800",
   304 => x"03060c18",
   305 => x"3060c000",
   306 => x"3c666e7e",
   307 => x"76663c00",
   308 => x"18387818",
   309 => x"18181800",
   310 => x"3c66060c",
   311 => x"18307e00",
   312 => x"3c66061c",
   313 => x"06663c00",
   314 => x"1c3c6ccc",
   315 => x"fe0c0c00",
   316 => x"7e607c06",
   317 => x"06663c00",
   318 => x"1c30607c",
   319 => x"66663c00",
   320 => x"7e06060c",
   321 => x"18181800",
   322 => x"3c66663c",
   323 => x"66663c00",
   324 => x"3c66663e",
   325 => x"060c3800",
   326 => x"00181800",
   327 => x"00181800",
   328 => x"00181800",
   329 => x"00181830",
   330 => x"00061860",
   331 => x"18060000",
   332 => x"00007e00",
   333 => x"7e000000",
   334 => x"00601806",
   335 => x"18600000",
   336 => x"3c66060c",
   337 => x"18001800",
   338 => x"7cc6ded6",
   339 => x"dec07800",
   340 => x"3c66667e",
   341 => x"66666600",
   342 => x"7c66667c",
   343 => x"66667c00",
   344 => x"1e306060",
   345 => x"60301e00",
   346 => x"786c6666",
   347 => x"666c7800",
   348 => x"7e606078",
   349 => x"60607e00",
   350 => x"7e606078",
   351 => x"60606000",
   352 => x"3c66606e",
   353 => x"66663e00",
   354 => x"6666667e",
   355 => x"66666600",
   356 => x"3c181818",
   357 => x"18183c00",
   358 => x"06060606",
   359 => x"06663c00",
   360 => x"c6ccd8f0",
   361 => x"d8ccc600",
   362 => x"60606060",
   363 => x"60607e00",
   364 => x"c6eefed6",
   365 => x"c6c6c600",
   366 => x"c6e6f6de",
   367 => x"cec6c600",
   368 => x"3c666666",
   369 => x"66663c00",
   370 => x"7c66667c",
   371 => x"60606000",
   372 => x"78cccccc",
   373 => x"ccdc7e00",
   374 => x"7c66667c",
   375 => x"6c666600",
   376 => x"3c66703c",
   377 => x"0e663c00",
   378 => x"7e181818",
   379 => x"18181800",
   380 => x"66666666",
   381 => x"66663c00",
   382 => x"66666666",
   383 => x"3c3c1800",
   384 => x"c6c6c6d6",
   385 => x"feeec600",
   386 => x"c3663c18",
   387 => x"3c66c300",
   388 => x"c3663c18",
   389 => x"18181800",
   390 => x"fe0c1830",
   391 => x"60c0fe00",
   392 => x"3c303030",
   393 => x"30303c00",
   394 => x"c0603018",
   395 => x"0c060300",
   396 => x"3c0c0c0c",
   397 => x"0c0c3c00",
   398 => x"10386cc6",
   399 => x"00000000",
   400 => x"00000000",
   401 => x"000000fe",
   402 => x"18180c00",
   403 => x"00000000",
   404 => x"00003c06",
   405 => x"3e663e00",
   406 => x"60607c66",
   407 => x"66667c00",
   408 => x"00003c60",
   409 => x"60603c00",
   410 => x"06063e66",
   411 => x"66663e00",
   412 => x"00003c66",
   413 => x"7e603c00",
   414 => x"1c307c30",
   415 => x"30303000",
   416 => x"00003e66",
   417 => x"663e063c",
   418 => x"60607c66",
   419 => x"66666600",
   420 => x"18001818",
   421 => x"18180c00",
   422 => x"0c000c0c",
   423 => x"0c0c0c78",
   424 => x"6060666c",
   425 => x"786c6600",
   426 => x"18181818",
   427 => x"18180c00",
   428 => x"0000ecfe",
   429 => x"d6c6c600",
   430 => x"00007c66",
   431 => x"66666600",
   432 => x"00003c66",
   433 => x"66663c00",
   434 => x"00007c66",
   435 => x"667c6060",
   436 => x"00003e66",
   437 => x"663e0606",
   438 => x"00007c66",
   439 => x"60606000",
   440 => x"00003c60",
   441 => x"3c067c00",
   442 => x"30307c30",
   443 => x"30301c00",
   444 => x"00006666",
   445 => x"66663e00",
   446 => x"00006666",
   447 => x"663c1800",
   448 => x"0000c6c6",
   449 => x"d6fe6c00",
   450 => x"0000c66c",
   451 => x"386cc600",
   452 => x"00006666",
   453 => x"663c1830",
   454 => x"00007e0c",
   455 => x"18307e00",
   456 => x"0e181870",
   457 => x"18180e00",
   458 => x"18181818",
   459 => x"18181800",
   460 => x"7018180e",
   461 => x"18187000",
   462 => x"729c0000",
   463 => x"00000000",
   464 => x"fefefefe",
   465 => x"fefefe00",
   466 => x"00000000",
   467 => x"00000000",
   468 => x"00000000",
   469 => x"00000000",
   470 => x"00000000",
   471 => x"00000000",
   472 => x"00000000",
   473 => x"00000000",
   474 => x"00000000",
   475 => x"00000000",
   476 => x"00000000",
   477 => x"00000000",
   478 => x"00000000",
   479 => x"00000000",
   480 => x"00000000",
   481 => x"00000000",
   482 => x"00000000",
   483 => x"00000000",
   484 => x"00000000",
   485 => x"00000000",
   486 => x"00000000",
   487 => x"00000000",
   488 => x"00000000",
   489 => x"00000000",
   490 => x"00000000",
   491 => x"00000000",
   492 => x"00000000",
   493 => x"00000000",
   494 => x"00000000",
   495 => x"00000000",
   496 => x"00000000",
   497 => x"00000000",
   498 => x"00000000",
   499 => x"00000000",
   500 => x"00000000",
   501 => x"00000000",
   502 => x"00000000",
   503 => x"00000000",
   504 => x"00000000",
   505 => x"00000000",
   506 => x"00000000",
   507 => x"00000000",
   508 => x"00000000",
   509 => x"00000000",
   510 => x"00000000",
   511 => x"00000000",
   512 => x"00000000",
   513 => x"00000000",
   514 => x"00000000",
   515 => x"00000000",
   516 => x"00000000",
   517 => x"00000000",
   518 => x"00000000",
   519 => x"00000000",
   520 => x"00000000",
   521 => x"00000000",
   522 => x"00000000",
   523 => x"00000000",
   524 => x"00000000",
   525 => x"00000000",
   526 => x"00000000",
   527 => x"00000000",
   528 => x"00000000",
   529 => x"00000000",
   530 => x"00000000",
   531 => x"00000000",
   532 => x"00000000",
   533 => x"00000000",
   534 => x"00000000",
   535 => x"00000000",
   536 => x"00000000",
   537 => x"00000000",
   538 => x"00000000",
   539 => x"00000000",
   540 => x"00000000",
   541 => x"00000000",
   542 => x"00000000",
   543 => x"00000000",
   544 => x"00000000",
   545 => x"00000000",
   546 => x"00000000",
   547 => x"00000000",
   548 => x"00000000",
   549 => x"00000000",
   550 => x"00000000",
   551 => x"00000000",
   552 => x"00000000",
   553 => x"00000000",
   554 => x"00000000",
   555 => x"00000000",
   556 => x"00000000",
   557 => x"00000000",
   558 => x"00000000",
   559 => x"00000000",
   560 => x"00000000",
   561 => x"00000000",
   562 => x"00000000",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

