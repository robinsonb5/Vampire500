-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"f2040000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"8cb07383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040ba0",
    29 => x"8080fd0b",
    30 => x"a0808ba6",
    31 => x"040ba080",
    32 => x"80fd0402",
    33 => x"f8050d73",
    34 => x"52ff8408",
    35 => x"70882a70",
    36 => x"81065151",
    37 => x"5170802e",
    38 => x"f03871ff",
    39 => x"840c71a0",
    40 => x"8092bc0c",
    41 => x"0288050d",
    42 => x"0402f005",
    43 => x"0d755380",
    44 => x"73a08080",
    45 => x"b42d7081",
    46 => x"ff065353",
    47 => x"5470742e",
    48 => x"b0387181",
    49 => x"ff068114",
    50 => x"5452ff84",
    51 => x"0870882a",
    52 => x"70810651",
    53 => x"51517080",
    54 => x"2ef03871",
    55 => x"ff840c81",
    56 => x"1473a080",
    57 => x"80b42d70",
    58 => x"81ff0653",
    59 => x"535470d2",
    60 => x"3873a080",
    61 => x"92bc0c02",
    62 => x"90050d04",
    63 => x"02c4050d",
    64 => x"0280c005",
    65 => x"a080939c",
    66 => x"5b568076",
    67 => x"70840558",
    68 => x"08715e5e",
    69 => x"577c7084",
    70 => x"055e0858",
    71 => x"805b7798",
    72 => x"2a78882b",
    73 => x"59537288",
    74 => x"38765ea0",
    75 => x"8084a504",
    76 => x"7b802e81",
    77 => x"ca38805c",
    78 => x"7280e42e",
    79 => x"9f387280",
    80 => x"e4268d38",
    81 => x"7280e32e",
    82 => x"80ee38a0",
    83 => x"8083c504",
    84 => x"7280f32e",
    85 => x"80cc38a0",
    86 => x"8083c504",
    87 => x"75841771",
    88 => x"087e5c56",
    89 => x"57528755",
    90 => x"739c2a74",
    91 => x"842b5552",
    92 => x"71802e83",
    93 => x"38815989",
    94 => x"72258938",
    95 => x"b71252a0",
    96 => x"80838704",
    97 => x"b0125278",
    98 => x"802e8838",
    99 => x"7151a080",
   100 => x"81832dff",
   101 => x"15557480",
   102 => x"25ce3880",
   103 => x"54a08083",
   104 => x"db047584",
   105 => x"17710870",
   106 => x"545c5752",
   107 => x"a08081a9",
   108 => x"2d7b54a0",
   109 => x"8083db04",
   110 => x"75841771",
   111 => x"08555752",
   112 => x"a080848e",
   113 => x"04a551a0",
   114 => x"8081832d",
   115 => x"7251a080",
   116 => x"81832d82",
   117 => x"1757a080",
   118 => x"84980473",
   119 => x"ff155552",
   120 => x"807225b4",
   121 => x"38797081",
   122 => x"055ba080",
   123 => x"80b42d70",
   124 => x"5253a080",
   125 => x"81832d81",
   126 => x"1757a080",
   127 => x"83db0472",
   128 => x"a52e0981",
   129 => x"06883881",
   130 => x"5ca08084",
   131 => x"98047251",
   132 => x"a0808183",
   133 => x"2d811757",
   134 => x"811b5b83",
   135 => x"7b25fdfe",
   136 => x"3872fdf1",
   137 => x"387da080",
   138 => x"92bc0c02",
   139 => x"bc050d04",
   140 => x"02f4050d",
   141 => x"74765253",
   142 => x"80712590",
   143 => x"38705272",
   144 => x"70840554",
   145 => x"08ff1353",
   146 => x"5171f438",
   147 => x"028c050d",
   148 => x"0402d805",
   149 => x"0d7b7d5b",
   150 => x"56810ba0",
   151 => x"808cc059",
   152 => x"57835977",
   153 => x"08760c75",
   154 => x"08780856",
   155 => x"5473752e",
   156 => x"92387508",
   157 => x"537452a0",
   158 => x"808cd051",
   159 => x"a08081fc",
   160 => x"2d805779",
   161 => x"527551a0",
   162 => x"8084b02d",
   163 => x"75085473",
   164 => x"752e9238",
   165 => x"75085374",
   166 => x"52a0808d",
   167 => x"9051a080",
   168 => x"81fc2d80",
   169 => x"57ff1984",
   170 => x"19595978",
   171 => x"8025ffb3",
   172 => x"3876a080",
   173 => x"92bc0c02",
   174 => x"a8050d04",
   175 => x"02ec050d",
   176 => x"76548155",
   177 => x"85aad5aa",
   178 => x"d5740cfa",
   179 => x"d5aad5aa",
   180 => x"0b8c150c",
   181 => x"cc74a080",
   182 => x"80c92db3",
   183 => x"0b8f15a0",
   184 => x"8080c92d",
   185 => x"73085372",
   186 => x"fce2d5aa",
   187 => x"d52e9038",
   188 => x"730852a0",
   189 => x"808dd051",
   190 => x"a08081fc",
   191 => x"2d80558c",
   192 => x"14085372",
   193 => x"fad5aad4",
   194 => x"b32e9138",
   195 => x"8c140852",
   196 => x"a0808e8c",
   197 => x"51a08081",
   198 => x"fc2d8055",
   199 => x"77527351",
   200 => x"a08084b0",
   201 => x"2d730853",
   202 => x"72fce2d5",
   203 => x"aad52e90",
   204 => x"38730852",
   205 => x"a0808ec8",
   206 => x"51a08081",
   207 => x"fc2d8055",
   208 => x"8c140853",
   209 => x"72fad5aa",
   210 => x"d4b32e91",
   211 => x"388c1408",
   212 => x"52a0808f",
   213 => x"8451a080",
   214 => x"81fc2d80",
   215 => x"5574a080",
   216 => x"92bc0c02",
   217 => x"94050d04",
   218 => x"02c4050d",
   219 => x"605e8062",
   220 => x"90808029",
   221 => x"ff05a080",
   222 => x"8fc0535e",
   223 => x"5ca08081",
   224 => x"fc2d80e1",
   225 => x"b35780fe",
   226 => x"5bae51a0",
   227 => x"8081832d",
   228 => x"76107096",
   229 => x"2a708106",
   230 => x"51565774",
   231 => x"802e8538",
   232 => x"76810757",
   233 => x"76952a70",
   234 => x"81065155",
   235 => x"74802e85",
   236 => x"38768132",
   237 => x"57787707",
   238 => x"7d06775b",
   239 => x"598fffff",
   240 => x"5876bfff",
   241 => x"ff06707a",
   242 => x"32822b7f",
   243 => x"11515776",
   244 => x"0c761070",
   245 => x"962a7081",
   246 => x"06515657",
   247 => x"74802e85",
   248 => x"38768107",
   249 => x"5776952a",
   250 => x"70810651",
   251 => x"5574802e",
   252 => x"85387681",
   253 => x"3257ff18",
   254 => x"58778025",
   255 => x"c4387957",
   256 => x"8fffff58",
   257 => x"76bfffff",
   258 => x"06707a32",
   259 => x"822b7f11",
   260 => x"70085151",
   261 => x"56567476",
   262 => x"2ea63880",
   263 => x"7c53a080",
   264 => x"8fd0525f",
   265 => x"a08081fc",
   266 => x"2d745475",
   267 => x"537552a0",
   268 => x"808fe451",
   269 => x"a08081fc",
   270 => x"2d7e5ca0",
   271 => x"8088c304",
   272 => x"811c5c76",
   273 => x"1070962a",
   274 => x"70810651",
   275 => x"56577480",
   276 => x"2e853876",
   277 => x"81075776",
   278 => x"952a7081",
   279 => x"06515574",
   280 => x"802e8538",
   281 => x"76813257",
   282 => x"ff185877",
   283 => x"8025ff94",
   284 => x"38ff1b5b",
   285 => x"7afe9238",
   286 => x"8a51a080",
   287 => x"81832d7e",
   288 => x"a08092bc",
   289 => x"0c02bc05",
   290 => x"0d0402d0",
   291 => x"050d7d5b",
   292 => x"815a8059",
   293 => x"80c07a59",
   294 => x"5c85ada9",
   295 => x"89bb7b0c",
   296 => x"79578156",
   297 => x"97557776",
   298 => x"07822b7b",
   299 => x"11515485",
   300 => x"ada989bb",
   301 => x"740c7510",
   302 => x"ff165656",
   303 => x"748025e6",
   304 => x"38771081",
   305 => x"18585898",
   306 => x"7725d738",
   307 => x"7e527a51",
   308 => x"a08084b0",
   309 => x"2d8158ff",
   310 => x"8787a5c3",
   311 => x"7b0c9757",
   312 => x"77822b7b",
   313 => x"11700856",
   314 => x"565673ff",
   315 => x"8787a5c3",
   316 => x"2e098106",
   317 => x"8a387878",
   318 => x"0759a080",
   319 => x"8a9c0474",
   320 => x"08547385",
   321 => x"ada989bb",
   322 => x"2e923880",
   323 => x"75085476",
   324 => x"53a08090",
   325 => x"8c525aa0",
   326 => x"8081fc2d",
   327 => x"7710ff18",
   328 => x"58587680",
   329 => x"25ffb938",
   330 => x"78822b59",
   331 => x"78802e80",
   332 => x"de387852",
   333 => x"a08090ac",
   334 => x"51a08081",
   335 => x"fc2d7899",
   336 => x"2a813270",
   337 => x"81067009",
   338 => x"81057072",
   339 => x"07700970",
   340 => x"9f2c7f06",
   341 => x"7e109fff",
   342 => x"fffe0662",
   343 => x"812a435f",
   344 => x"5f515156",
   345 => x"515578d6",
   346 => x"38790981",
   347 => x"05707b07",
   348 => x"9f2a5154",
   349 => x"7bbf2695",
   350 => x"3873802e",
   351 => x"9038a080",
   352 => x"90c451a0",
   353 => x"8081fc2d",
   354 => x"a0808b8f",
   355 => x"04815c7b",
   356 => x"52a08091",
   357 => x"9051a080",
   358 => x"81fc2d7b",
   359 => x"a08092bc",
   360 => x"0c02b005",
   361 => x"0d0402f4",
   362 => x"050d88bd",
   363 => x"0bff880c",
   364 => x"a0805280",
   365 => x"51a08084",
   366 => x"d12da080",
   367 => x"92bc0880",
   368 => x"2e8b38a0",
   369 => x"8091cc51",
   370 => x"a08081fc",
   371 => x"2da08052",
   372 => x"8051a080",
   373 => x"85bc2da0",
   374 => x"8092bc08",
   375 => x"802e8b38",
   376 => x"a08091f0",
   377 => x"51a08081",
   378 => x"fc2da080",
   379 => x"528051a0",
   380 => x"80898a2d",
   381 => x"a08092bc",
   382 => x"0853a080",
   383 => x"92bc0880",
   384 => x"2e8b38a0",
   385 => x"80928c51",
   386 => x"a08081fc",
   387 => x"2d725280",
   388 => x"51a08086",
   389 => x"e82da080",
   390 => x"92bc0880",
   391 => x"2eff9138",
   392 => x"a08092a4",
   393 => x"51a08081",
   394 => x"fc2da080",
   395 => x"8bb00400",
   396 => x"00ffffff",
   397 => x"ff00ffff",
   398 => x"ffff00ff",
   399 => x"ffffff00",
   400 => x"00000000",
   401 => x"55555555",
   402 => x"aaaaaaaa",
   403 => x"ffffffff",
   404 => x"53616e69",
   405 => x"74792063",
   406 => x"6865636b",
   407 => x"20666169",
   408 => x"6c656420",
   409 => x"28626566",
   410 => x"6f726520",
   411 => x"63616368",
   412 => x"65207265",
   413 => x"66726573",
   414 => x"6829206f",
   415 => x"6e203078",
   416 => x"25642028",
   417 => x"676f7420",
   418 => x"30782564",
   419 => x"290a0000",
   420 => x"53616e69",
   421 => x"74792063",
   422 => x"6865636b",
   423 => x"20666169",
   424 => x"6c656420",
   425 => x"28616674",
   426 => x"65722063",
   427 => x"61636865",
   428 => x"20726566",
   429 => x"72657368",
   430 => x"29206f6e",
   431 => x"20307825",
   432 => x"64202867",
   433 => x"6f742030",
   434 => x"78256429",
   435 => x"0a000000",
   436 => x"42797465",
   437 => x"20636865",
   438 => x"636b2066",
   439 => x"61696c65",
   440 => x"64202862",
   441 => x"65666f72",
   442 => x"65206361",
   443 => x"63686520",
   444 => x"72656672",
   445 => x"65736829",
   446 => x"20617420",
   447 => x"30202867",
   448 => x"6f742030",
   449 => x"78256429",
   450 => x"0a000000",
   451 => x"42797465",
   452 => x"20636865",
   453 => x"636b2066",
   454 => x"61696c65",
   455 => x"64202862",
   456 => x"65666f72",
   457 => x"65206361",
   458 => x"63686520",
   459 => x"72656672",
   460 => x"65736829",
   461 => x"20617420",
   462 => x"33202867",
   463 => x"6f742030",
   464 => x"78256429",
   465 => x"0a000000",
   466 => x"42797465",
   467 => x"20636865",
   468 => x"636b2066",
   469 => x"61696c65",
   470 => x"64202861",
   471 => x"66746572",
   472 => x"20636163",
   473 => x"68652072",
   474 => x"65667265",
   475 => x"73682920",
   476 => x"61742030",
   477 => x"2028676f",
   478 => x"74203078",
   479 => x"2564290a",
   480 => x"00000000",
   481 => x"42797465",
   482 => x"20636865",
   483 => x"636b2066",
   484 => x"61696c65",
   485 => x"64202861",
   486 => x"66746572",
   487 => x"20636163",
   488 => x"68652072",
   489 => x"65667265",
   490 => x"73682920",
   491 => x"61742033",
   492 => x"2028676f",
   493 => x"74203078",
   494 => x"2564290a",
   495 => x"00000000",
   496 => x"43686563",
   497 => x"6b696e67",
   498 => x"206d656d",
   499 => x"6f727900",
   500 => x"30782564",
   501 => x"20676f6f",
   502 => x"64207265",
   503 => x"6164732c",
   504 => x"20000000",
   505 => x"4572726f",
   506 => x"72206174",
   507 => x"20307825",
   508 => x"642c2065",
   509 => x"78706563",
   510 => x"74656420",
   511 => x"30782564",
   512 => x"2c20676f",
   513 => x"74203078",
   514 => x"25640a00",
   515 => x"42616420",
   516 => x"64617461",
   517 => x"20666f75",
   518 => x"6e642061",
   519 => x"74203078",
   520 => x"25642028",
   521 => x"30782564",
   522 => x"290a0000",
   523 => x"416c6961",
   524 => x"73657320",
   525 => x"666f756e",
   526 => x"64206174",
   527 => x"20307825",
   528 => x"640a0000",
   529 => x"28416c69",
   530 => x"61736573",
   531 => x"2070726f",
   532 => x"6261626c",
   533 => x"79207369",
   534 => x"6d706c79",
   535 => x"20696e64",
   536 => x"69636174",
   537 => x"65207468",
   538 => x"61742052",
   539 => x"414d0a69",
   540 => x"7320736d",
   541 => x"616c6c65",
   542 => x"72207468",
   543 => x"616e2036",
   544 => x"34206d65",
   545 => x"67616279",
   546 => x"74657329",
   547 => x"0a000000",
   548 => x"53445241",
   549 => x"4d207369",
   550 => x"7a652028",
   551 => x"61737375",
   552 => x"6d696e67",
   553 => x"206e6f20",
   554 => x"61646472",
   555 => x"65737320",
   556 => x"6661756c",
   557 => x"74732920",
   558 => x"69732030",
   559 => x"78256420",
   560 => x"6d656761",
   561 => x"62797465",
   562 => x"730a0000",
   563 => x"46697273",
   564 => x"74207374",
   565 => x"61676520",
   566 => x"73616e69",
   567 => x"74792063",
   568 => x"6865636b",
   569 => x"20706173",
   570 => x"7365642e",
   571 => x"0a000000",
   572 => x"42797465",
   573 => x"20286471",
   574 => x"6d292063",
   575 => x"6865636b",
   576 => x"20706173",
   577 => x"7365640a",
   578 => x"00000000",
   579 => x"41646472",
   580 => x"65737320",
   581 => x"63686563",
   582 => x"6b207061",
   583 => x"73736564",
   584 => x"2e0a0000",
   585 => x"4c465352",
   586 => x"20636865",
   587 => x"636b2070",
   588 => x"61737365",
   589 => x"642e0a0a",
   590 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

