library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package sdram_config is

constant sdram_rows : integer := 13;
constant sdram_cols : integer := 9;

end package;
