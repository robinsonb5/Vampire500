-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"f2040000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"8cf87383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040ba0",
    29 => x"8080fd0b",
    30 => x"a0808beb",
    31 => x"040ba080",
    32 => x"80fd0402",
    33 => x"f8050d73",
    34 => x"52ff8408",
    35 => x"70882a70",
    36 => x"81065151",
    37 => x"5170802e",
    38 => x"f03871ff",
    39 => x"840c71a0",
    40 => x"8093840c",
    41 => x"0288050d",
    42 => x"0402f005",
    43 => x"0d755380",
    44 => x"73a08080",
    45 => x"b42d7081",
    46 => x"ff065353",
    47 => x"5470742e",
    48 => x"b0387181",
    49 => x"ff068114",
    50 => x"5452ff84",
    51 => x"0870882a",
    52 => x"70810651",
    53 => x"51517080",
    54 => x"2ef03871",
    55 => x"ff840c81",
    56 => x"1473a080",
    57 => x"80b42d70",
    58 => x"81ff0653",
    59 => x"535470d2",
    60 => x"3873a080",
    61 => x"93840c02",
    62 => x"90050d04",
    63 => x"02c4050d",
    64 => x"0280c005",
    65 => x"a08093e4",
    66 => x"5b568076",
    67 => x"70840558",
    68 => x"08715e5e",
    69 => x"577c7084",
    70 => x"055e0858",
    71 => x"805b7798",
    72 => x"2a78882b",
    73 => x"59537288",
    74 => x"38765ea0",
    75 => x"8084a504",
    76 => x"7b802e81",
    77 => x"ca38805c",
    78 => x"7280e42e",
    79 => x"9f387280",
    80 => x"e4268d38",
    81 => x"7280e32e",
    82 => x"80ee38a0",
    83 => x"8083c504",
    84 => x"7280f32e",
    85 => x"80cc38a0",
    86 => x"8083c504",
    87 => x"75841771",
    88 => x"087e5c56",
    89 => x"57528755",
    90 => x"739c2a74",
    91 => x"842b5552",
    92 => x"71802e83",
    93 => x"38815989",
    94 => x"72258938",
    95 => x"b71252a0",
    96 => x"80838704",
    97 => x"b0125278",
    98 => x"802e8838",
    99 => x"7151a080",
   100 => x"81832dff",
   101 => x"15557480",
   102 => x"25ce3880",
   103 => x"54a08083",
   104 => x"db047584",
   105 => x"17710870",
   106 => x"545c5752",
   107 => x"a08081a9",
   108 => x"2d7b54a0",
   109 => x"8083db04",
   110 => x"75841771",
   111 => x"08555752",
   112 => x"a080848e",
   113 => x"04a551a0",
   114 => x"8081832d",
   115 => x"7251a080",
   116 => x"81832d82",
   117 => x"1757a080",
   118 => x"84980473",
   119 => x"ff155552",
   120 => x"807225b4",
   121 => x"38797081",
   122 => x"055ba080",
   123 => x"80b42d70",
   124 => x"5253a080",
   125 => x"81832d81",
   126 => x"1757a080",
   127 => x"83db0472",
   128 => x"a52e0981",
   129 => x"06883881",
   130 => x"5ca08084",
   131 => x"98047251",
   132 => x"a0808183",
   133 => x"2d811757",
   134 => x"811b5b83",
   135 => x"7b25fdfe",
   136 => x"3872fdf1",
   137 => x"387da080",
   138 => x"93840c02",
   139 => x"bc050d04",
   140 => x"02f4050d",
   141 => x"74765253",
   142 => x"80712590",
   143 => x"38705272",
   144 => x"70840554",
   145 => x"08ff1353",
   146 => x"5171f438",
   147 => x"028c050d",
   148 => x"0402d805",
   149 => x"0d7b7d5b",
   150 => x"56810ba0",
   151 => x"808d8859",
   152 => x"57835977",
   153 => x"08760c75",
   154 => x"08780856",
   155 => x"5473752e",
   156 => x"92387508",
   157 => x"537452a0",
   158 => x"808d9851",
   159 => x"a08081fc",
   160 => x"2d805779",
   161 => x"527551a0",
   162 => x"8084b02d",
   163 => x"75085473",
   164 => x"752e9238",
   165 => x"75085374",
   166 => x"52a0808d",
   167 => x"d851a080",
   168 => x"81fc2d80",
   169 => x"57ff1984",
   170 => x"19595978",
   171 => x"8025ffb3",
   172 => x"3876a080",
   173 => x"93840c02",
   174 => x"a8050d04",
   175 => x"02ec050d",
   176 => x"76548155",
   177 => x"85aad5aa",
   178 => x"d5740cfa",
   179 => x"d5aad5aa",
   180 => x"0b8c150c",
   181 => x"cc74a080",
   182 => x"80c92db3",
   183 => x"0b8f15a0",
   184 => x"8080c92d",
   185 => x"73085372",
   186 => x"fce2d5aa",
   187 => x"d52e9038",
   188 => x"730852a0",
   189 => x"808e9851",
   190 => x"a08081fc",
   191 => x"2d80558c",
   192 => x"14085372",
   193 => x"fad5aad4",
   194 => x"b32e9138",
   195 => x"8c140852",
   196 => x"a0808ed4",
   197 => x"51a08081",
   198 => x"fc2d8055",
   199 => x"77527351",
   200 => x"a08084b0",
   201 => x"2d730853",
   202 => x"72fce2d5",
   203 => x"aad52e90",
   204 => x"38730852",
   205 => x"a0808f90",
   206 => x"51a08081",
   207 => x"fc2d8055",
   208 => x"8c140853",
   209 => x"72fad5aa",
   210 => x"d4b32e91",
   211 => x"388c1408",
   212 => x"52a0808f",
   213 => x"cc51a080",
   214 => x"81fc2d80",
   215 => x"5574a080",
   216 => x"93840c02",
   217 => x"94050d04",
   218 => x"02c8050d",
   219 => x"7f5c800b",
   220 => x"a0809088",
   221 => x"525ba080",
   222 => x"81fc2d80",
   223 => x"e1b3578e",
   224 => x"5d76598f",
   225 => x"ffff5a76",
   226 => x"bfffff06",
   227 => x"77107096",
   228 => x"2a708106",
   229 => x"51575858",
   230 => x"74802e85",
   231 => x"38768107",
   232 => x"5776952a",
   233 => x"70810651",
   234 => x"5574802e",
   235 => x"85387681",
   236 => x"325776bf",
   237 => x"ffff0678",
   238 => x"84291d79",
   239 => x"710c5670",
   240 => x"84291d56",
   241 => x"750c7610",
   242 => x"70962a70",
   243 => x"81065156",
   244 => x"5774802e",
   245 => x"85387681",
   246 => x"07577695",
   247 => x"2a708106",
   248 => x"51557480",
   249 => x"2e853876",
   250 => x"813257ff",
   251 => x"1a5a7980",
   252 => x"25ff9438",
   253 => x"78578fff",
   254 => x"ff5a76bf",
   255 => x"ffff0677",
   256 => x"1070962a",
   257 => x"70810651",
   258 => x"57585674",
   259 => x"802e8538",
   260 => x"76810757",
   261 => x"76952a70",
   262 => x"81065155",
   263 => x"74802e85",
   264 => x"38768132",
   265 => x"5776bfff",
   266 => x"ff067684",
   267 => x"291d7008",
   268 => x"575a5874",
   269 => x"762ea738",
   270 => x"807b53a0",
   271 => x"80909c52",
   272 => x"5ea08081",
   273 => x"fc2d7808",
   274 => x"54755375",
   275 => x"52a08090",
   276 => x"b051a080",
   277 => x"81fc2d7d",
   278 => x"5ba08088",
   279 => x"e104811b",
   280 => x"5b778429",
   281 => x"1c700856",
   282 => x"5674782e",
   283 => x"a738807b",
   284 => x"53a08090",
   285 => x"9c525ea0",
   286 => x"8081fc2d",
   287 => x"75085477",
   288 => x"537752a0",
   289 => x"8090b051",
   290 => x"a08081fc",
   291 => x"2d7d5ba0",
   292 => x"80899704",
   293 => x"811b5b76",
   294 => x"1070962a",
   295 => x"70810651",
   296 => x"56577480",
   297 => x"2e853876",
   298 => x"81075776",
   299 => x"952a7081",
   300 => x"06515574",
   301 => x"802e8538",
   302 => x"76813257",
   303 => x"ff1a5a79",
   304 => x"8025feb6",
   305 => x"38ff1d5d",
   306 => x"7cfdb638",
   307 => x"7da08093",
   308 => x"840c02b8",
   309 => x"050d0402",
   310 => x"cc050d7e",
   311 => x"5c815b80",
   312 => x"5a80c07b",
   313 => x"585d85ad",
   314 => x"a989bb7c",
   315 => x"0c7a5681",
   316 => x"58975576",
   317 => x"7807822b",
   318 => x"7c115154",
   319 => x"85ada989",
   320 => x"bb740c77",
   321 => x"10ff1656",
   322 => x"58748025",
   323 => x"e6387610",
   324 => x"81175757",
   325 => x"987625d7",
   326 => x"387f527b",
   327 => x"51a08084",
   328 => x"b02d8157",
   329 => x"ff8787a5",
   330 => x"c37c0c97",
   331 => x"56807782",
   332 => x"2b7d1170",
   333 => x"0857575a",
   334 => x"5873ff87",
   335 => x"87a5c32e",
   336 => x"0981068a",
   337 => x"38797707",
   338 => x"5aa0808a",
   339 => x"eb047408",
   340 => x"547385ad",
   341 => x"a989bb2e",
   342 => x"92387775",
   343 => x"08547953",
   344 => x"a08090d8",
   345 => x"525ba080",
   346 => x"81fc2d76",
   347 => x"10ff1757",
   348 => x"57758025",
   349 => x"ffb73879",
   350 => x"802eba38",
   351 => x"79822b52",
   352 => x"a08090f8",
   353 => x"51a08081",
   354 => x"fc2d7999",
   355 => x"2a813270",
   356 => x"81067009",
   357 => x"81057072",
   358 => x"07700970",
   359 => x"9f2c6006",
   360 => x"7f1087ff",
   361 => x"fffe0663",
   362 => x"812c4440",
   363 => x"40515156",
   364 => x"515579d6",
   365 => x"387a0981",
   366 => x"05707c07",
   367 => x"9f2a5154",
   368 => x"7cbf2490",
   369 => x"3873802e",
   370 => x"8b38a080",
   371 => x"919051a0",
   372 => x"8081fc2d",
   373 => x"7c52a080",
   374 => x"91dc51a0",
   375 => x"8081fc2d",
   376 => x"7aa08093",
   377 => x"840c02b4",
   378 => x"050d0402",
   379 => x"f8050d88",
   380 => x"bd0bff88",
   381 => x"0ca08052",
   382 => x"8051a080",
   383 => x"84d12da0",
   384 => x"80938408",
   385 => x"802e8b38",
   386 => x"a0809298",
   387 => x"51a08081",
   388 => x"fc2da080",
   389 => x"528051a0",
   390 => x"8085bc2d",
   391 => x"a0809384",
   392 => x"08802e8b",
   393 => x"38a08092",
   394 => x"bc51a080",
   395 => x"81fc2da0",
   396 => x"80528051",
   397 => x"a08089d7",
   398 => x"2da08093",
   399 => x"8408802e",
   400 => x"8b38a080",
   401 => x"92d851a0",
   402 => x"8081fc2d",
   403 => x"8051a080",
   404 => x"86e82da0",
   405 => x"80938408",
   406 => x"802e8b38",
   407 => x"a08092f0",
   408 => x"51a08081",
   409 => x"fc2da080",
   410 => x"8ed051a0",
   411 => x"8081fc2d",
   412 => x"a0808bf5",
   413 => x"04000000",
   414 => x"00ffffff",
   415 => x"ff00ffff",
   416 => x"ffff00ff",
   417 => x"ffffff00",
   418 => x"00000000",
   419 => x"55555555",
   420 => x"aaaaaaaa",
   421 => x"ffffffff",
   422 => x"53616e69",
   423 => x"74792063",
   424 => x"6865636b",
   425 => x"20666169",
   426 => x"6c656420",
   427 => x"28626566",
   428 => x"6f726520",
   429 => x"63616368",
   430 => x"65207265",
   431 => x"66726573",
   432 => x"6829206f",
   433 => x"6e203078",
   434 => x"25642028",
   435 => x"676f7420",
   436 => x"30782564",
   437 => x"290a0000",
   438 => x"53616e69",
   439 => x"74792063",
   440 => x"6865636b",
   441 => x"20666169",
   442 => x"6c656420",
   443 => x"28616674",
   444 => x"65722063",
   445 => x"61636865",
   446 => x"20726566",
   447 => x"72657368",
   448 => x"29206f6e",
   449 => x"20307825",
   450 => x"64202867",
   451 => x"6f742030",
   452 => x"78256429",
   453 => x"0a000000",
   454 => x"42797465",
   455 => x"20636865",
   456 => x"636b2066",
   457 => x"61696c65",
   458 => x"64202862",
   459 => x"65666f72",
   460 => x"65206361",
   461 => x"63686520",
   462 => x"72656672",
   463 => x"65736829",
   464 => x"20617420",
   465 => x"30202867",
   466 => x"6f742030",
   467 => x"78256429",
   468 => x"0a000000",
   469 => x"42797465",
   470 => x"20636865",
   471 => x"636b2066",
   472 => x"61696c65",
   473 => x"64202862",
   474 => x"65666f72",
   475 => x"65206361",
   476 => x"63686520",
   477 => x"72656672",
   478 => x"65736829",
   479 => x"20617420",
   480 => x"33202867",
   481 => x"6f742030",
   482 => x"78256429",
   483 => x"0a000000",
   484 => x"42797465",
   485 => x"20636865",
   486 => x"636b2066",
   487 => x"61696c65",
   488 => x"64202861",
   489 => x"66746572",
   490 => x"20636163",
   491 => x"68652072",
   492 => x"65667265",
   493 => x"73682920",
   494 => x"61742030",
   495 => x"2028676f",
   496 => x"74203078",
   497 => x"2564290a",
   498 => x"00000000",
   499 => x"42797465",
   500 => x"20636865",
   501 => x"636b2066",
   502 => x"61696c65",
   503 => x"64202861",
   504 => x"66746572",
   505 => x"20636163",
   506 => x"68652072",
   507 => x"65667265",
   508 => x"73682920",
   509 => x"61742033",
   510 => x"2028676f",
   511 => x"74203078",
   512 => x"2564290a",
   513 => x"00000000",
   514 => x"43686563",
   515 => x"6b696e67",
   516 => x"206d656d",
   517 => x"6f72792e",
   518 => x"2e2e0a00",
   519 => x"30782564",
   520 => x"20676f6f",
   521 => x"64207265",
   522 => x"6164732c",
   523 => x"20000000",
   524 => x"4572726f",
   525 => x"72206174",
   526 => x"20307825",
   527 => x"642c2065",
   528 => x"78706563",
   529 => x"74656420",
   530 => x"30782564",
   531 => x"2c20676f",
   532 => x"74203078",
   533 => x"25640a00",
   534 => x"42616420",
   535 => x"64617461",
   536 => x"20666f75",
   537 => x"6e642061",
   538 => x"74203078",
   539 => x"25642028",
   540 => x"30782564",
   541 => x"290a0000",
   542 => x"416c6961",
   543 => x"73657320",
   544 => x"666f756e",
   545 => x"64206174",
   546 => x"20307825",
   547 => x"640a0000",
   548 => x"28416c69",
   549 => x"61736573",
   550 => x"2070726f",
   551 => x"6261626c",
   552 => x"79207369",
   553 => x"6d706c79",
   554 => x"20696e64",
   555 => x"69636174",
   556 => x"65207468",
   557 => x"61742052",
   558 => x"414d2069",
   559 => x"7320736d",
   560 => x"616c6c65",
   561 => x"72207468",
   562 => x"616e2036",
   563 => x"34206d65",
   564 => x"67616279",
   565 => x"74657329",
   566 => x"00000000",
   567 => x"53445241",
   568 => x"4d207369",
   569 => x"7a652028",
   570 => x"61737375",
   571 => x"6d696e67",
   572 => x"206e6f20",
   573 => x"61646472",
   574 => x"65737320",
   575 => x"6661756c",
   576 => x"74732920",
   577 => x"69732030",
   578 => x"78256420",
   579 => x"6d656761",
   580 => x"62797465",
   581 => x"730a0000",
   582 => x"46697273",
   583 => x"74207374",
   584 => x"61676520",
   585 => x"73616e69",
   586 => x"74792063",
   587 => x"6865636b",
   588 => x"20706173",
   589 => x"7365642e",
   590 => x"0a000000",
   591 => x"42797465",
   592 => x"20286471",
   593 => x"6d292063",
   594 => x"6865636b",
   595 => x"20706173",
   596 => x"7365640a",
   597 => x"00000000",
   598 => x"41646472",
   599 => x"65737320",
   600 => x"63686563",
   601 => x"6b207061",
   602 => x"73736564",
   603 => x"2e0a0000",
   604 => x"4c465352",
   605 => x"20636865",
   606 => x"636b2070",
   607 => x"61737365",
   608 => x"642e0a00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

