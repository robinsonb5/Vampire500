-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08080f4",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"8bf87383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"800ba080",
    30 => x"8acc0c04",
    31 => x"ff3d0d83",
    32 => x"82800ba0",
    33 => x"808bb40c",
    34 => x"fea0800b",
    35 => x"86ffe280",
    36 => x"23800b86",
    37 => x"ffe28223",
    38 => x"800b86ff",
    39 => x"e2842380",
    40 => x"0b86ffe2",
    41 => x"8823800b",
    42 => x"86ffe28a",
    43 => x"23828080",
    44 => x"52a0bf51",
    45 => x"80727084",
    46 => x"05540cff",
    47 => x"11517080",
    48 => x"25f238bc",
    49 => x"0b86ffe1",
    50 => x"922381d4",
    51 => x"0b86ffe1",
    52 => x"942380d9",
    53 => x"810b86ff",
    54 => x"e18e23e9",
    55 => x"c10b86ff",
    56 => x"e1902386",
    57 => x"ff0b86ff",
    58 => x"e380239f",
    59 => x"ff0b86ff",
    60 => x"e38223a0",
    61 => x"808bb408",
    62 => x"70535181",
    63 => x"e0727082",
    64 => x"05542380",
    65 => x"72708205",
    66 => x"542381e2",
    67 => x"72708205",
    68 => x"5423fe80",
    69 => x"80727082",
    70 => x"055423ff",
    71 => x"72708205",
    72 => x"5423fe72",
    73 => x"2370902c",
    74 => x"527186ff",
    75 => x"e1802370",
    76 => x"86ffe182",
    77 => x"23800b86",
    78 => x"ffe18823",
    79 => x"fe87900b",
    80 => x"86ffe196",
    81 => x"23800ba0",
    82 => x"808adc0c",
    83 => x"800ba080",
    84 => x"8ae00c83",
    85 => x"3d0d04fb",
    86 => x"3d0d029f",
    87 => x"0533a080",
    88 => x"8ae008b1",
    89 => x"800a29a0",
    90 => x"808adc08",
    91 => x"0571a029",
    92 => x"16f88011",
    93 => x"08f88412",
    94 => x"08525757",
    95 => x"54567373",
    96 => x"3473ffb0",
    97 => x"143473fe",
    98 => x"e0143473",
    99 => x"fe901434",
   100 => x"74fdc014",
   101 => x"3474fcf0",
   102 => x"143474fc",
   103 => x"a0143474",
   104 => x"fbd01434",
   105 => x"758a2e80",
   106 => x"f138a080",
   107 => x"8adc0881",
   108 => x"05a0808a",
   109 => x"dc0ca080",
   110 => x"8adc0880",
   111 => x"d02eb838",
   112 => x"a0808ae0",
   113 => x"08992e85",
   114 => x"38873d0d",
   115 => x"04828080",
   116 => x"55828580",
   117 => x"549f9f53",
   118 => x"73708405",
   119 => x"55087570",
   120 => x"8405570c",
   121 => x"ff135372",
   122 => x"8025ed38",
   123 => x"980ba080",
   124 => x"8ae00c87",
   125 => x"3d0d04a0",
   126 => x"808ae008",
   127 => x"8105a080",
   128 => x"8ae00c80",
   129 => x"0ba0808a",
   130 => x"dc0ca080",
   131 => x"8ae00899",
   132 => x"2e098106",
   133 => x"ffb338ff",
   134 => x"b439a080",
   135 => x"8ae00881",
   136 => x"05a0808a",
   137 => x"e00ca080",
   138 => x"8ae00899",
   139 => x"2e098106",
   140 => x"ff9738ff",
   141 => x"9839f83d",
   142 => x"0d7a7070",
   143 => x"81055233",
   144 => x"58597680",
   145 => x"2e80fa38",
   146 => x"a0808ae0",
   147 => x"08b1800a",
   148 => x"29a0808a",
   149 => x"dc080577",
   150 => x"a02919f8",
   151 => x"801108f8",
   152 => x"84120859",
   153 => x"57f88805",
   154 => x"59547474",
   155 => x"3474ffb0",
   156 => x"153474fe",
   157 => x"e0153474",
   158 => x"fe901534",
   159 => x"75fdc015",
   160 => x"3475fcf0",
   161 => x"153475fc",
   162 => x"a0153475",
   163 => x"fbd01534",
   164 => x"768a2e81",
   165 => x"8238a080",
   166 => x"8adc0881",
   167 => x"05a0808a",
   168 => x"dc0ca080",
   169 => x"8adc0880",
   170 => x"d02e80c8",
   171 => x"38a0808a",
   172 => x"e008992e",
   173 => x"90387870",
   174 => x"81055a33",
   175 => x"5776ff88",
   176 => x"388a3d0d",
   177 => x"04828080",
   178 => x"55828580",
   179 => x"549f9f53",
   180 => x"73708405",
   181 => x"55087570",
   182 => x"8405570c",
   183 => x"ff135372",
   184 => x"8025ed38",
   185 => x"980ba080",
   186 => x"8ae00c78",
   187 => x"7081055a",
   188 => x"3357ca39",
   189 => x"a0808ae0",
   190 => x"088105a0",
   191 => x"808ae00c",
   192 => x"800ba080",
   193 => x"8adc0ca0",
   194 => x"808ae008",
   195 => x"992e0981",
   196 => x"06ffa338",
   197 => x"ffaf39a0",
   198 => x"808ae008",
   199 => x"8105a080",
   200 => x"8ae00ca0",
   201 => x"808ae008",
   202 => x"992e0981",
   203 => x"06ff8738",
   204 => x"ff9339ff",
   205 => x"3d0d028f",
   206 => x"053352ff",
   207 => x"84087088",
   208 => x"2a708106",
   209 => x"51515170",
   210 => x"802ef038",
   211 => x"71ff840c",
   212 => x"833d0d04",
   213 => x"fe3d0d74",
   214 => x"70335253",
   215 => x"70802ea1",
   216 => x"38705281",
   217 => x"1353ff84",
   218 => x"0870882a",
   219 => x"70810651",
   220 => x"51517080",
   221 => x"2ef03871",
   222 => x"ff840c72",
   223 => x"335271e3",
   224 => x"38843d0d",
   225 => x"04ff3d0d",
   226 => x"ff840870",
   227 => x"892a7081",
   228 => x"06515252",
   229 => x"70802ef0",
   230 => x"387181ff",
   231 => x"06a0808a",
   232 => x"cc0c833d",
   233 => x"0d04ff3d",
   234 => x"0d028f05",
   235 => x"3352ff84",
   236 => x"0870882a",
   237 => x"70810651",
   238 => x"51517080",
   239 => x"2ef03871",
   240 => x"ff840c83",
   241 => x"3d0d04f5",
   242 => x"3d0d8e3d",
   243 => x"70708405",
   244 => x"5208a080",
   245 => x"87a65b55",
   246 => x"5b807470",
   247 => x"81055633",
   248 => x"755a5457",
   249 => x"72772ebe",
   250 => x"3872a52e",
   251 => x"09810680",
   252 => x"c8387770",
   253 => x"81055933",
   254 => x"537280e4",
   255 => x"2e81b938",
   256 => x"7280e424",
   257 => x"80c93872",
   258 => x"80e32ea4",
   259 => x"388052a5",
   260 => x"51782d80",
   261 => x"52725178",
   262 => x"2d821757",
   263 => x"77708105",
   264 => x"59335372",
   265 => x"c43876a0",
   266 => x"808acc0c",
   267 => x"8d3d0d04",
   268 => x"7a841c83",
   269 => x"1233555c",
   270 => x"56805272",
   271 => x"51782d81",
   272 => x"17787081",
   273 => x"055a3354",
   274 => x"5772ff9d",
   275 => x"38d83972",
   276 => x"80f32e09",
   277 => x"8106ffb5",
   278 => x"387a841c",
   279 => x"7108585c",
   280 => x"54807633",
   281 => x"5b557975",
   282 => x"2e8d3881",
   283 => x"15701770",
   284 => x"33555b55",
   285 => x"72f538ff",
   286 => x"15548075",
   287 => x"25ff9d38",
   288 => x"75708105",
   289 => x"57335380",
   290 => x"52725178",
   291 => x"2d811774",
   292 => x"ff165656",
   293 => x"57807525",
   294 => x"ff823875",
   295 => x"70810557",
   296 => x"33538052",
   297 => x"7251782d",
   298 => x"811774ff",
   299 => x"16565657",
   300 => x"748024cc",
   301 => x"38fee539",
   302 => x"7a841c71",
   303 => x"08a0808b",
   304 => x"b80ba080",
   305 => x"8ae4545d",
   306 => x"565c5580",
   307 => x"5673762e",
   308 => x"098106bb",
   309 => x"38b00ba0",
   310 => x"808ae434",
   311 => x"811555ff",
   312 => x"15557433",
   313 => x"7a708105",
   314 => x"5c348116",
   315 => x"5674a080",
   316 => x"8ae42e09",
   317 => x"8106e838",
   318 => x"807a3475",
   319 => x"a0808bb8",
   320 => x"0bff1256",
   321 => x"57557480",
   322 => x"24fef538",
   323 => x"fe8e3973",
   324 => x"8f06a080",
   325 => x"9a880553",
   326 => x"72337570",
   327 => x"81055734",
   328 => x"73842a54",
   329 => x"73e93874",
   330 => x"a0808ae4",
   331 => x"2eca38ff",
   332 => x"15557433",
   333 => x"7a708105",
   334 => x"5c348116",
   335 => x"5674a080",
   336 => x"8ae42eff",
   337 => x"b338ff97",
   338 => x"39000000",
   339 => x"00000000",
   340 => x"00000000",
   341 => x"00000000",
   342 => x"00000000",
   343 => x"00000000",
   344 => x"00000000",
   345 => x"00000000",
   346 => x"00000000",
   347 => x"00000000",
   348 => x"00000000",
   349 => x"00000000",
   350 => x"00000000",
   351 => x"00000000",
   352 => x"00000000",
   353 => x"00000000",
   354 => x"00000000",
   355 => x"00000000",
   356 => x"00000000",
   357 => x"00000000",
   358 => x"00000000",
   359 => x"00000000",
   360 => x"00000000",
   361 => x"00000000",
   362 => x"00000000",
   363 => x"00000000",
   364 => x"00000000",
   365 => x"00000000",
   366 => x"00000000",
   367 => x"00000000",
   368 => x"00000000",
   369 => x"00000000",
   370 => x"00000000",
   371 => x"00000000",
   372 => x"00000000",
   373 => x"00000000",
   374 => x"00000000",
   375 => x"00000000",
   376 => x"00000000",
   377 => x"00000000",
   378 => x"00000000",
   379 => x"00000000",
   380 => x"00000000",
   381 => x"00000000",
   382 => x"00ffffff",
   383 => x"ff00ffff",
   384 => x"ffff00ff",
   385 => x"ffffff00",
   386 => x"00000000",
   387 => x"00000000",
   388 => x"18181818",
   389 => x"18001800",
   390 => x"6c6c0000",
   391 => x"00000000",
   392 => x"6c6cfe6c",
   393 => x"fe6c6c00",
   394 => x"183e603c",
   395 => x"067c1800",
   396 => x"0066acd8",
   397 => x"366acc00",
   398 => x"386c6876",
   399 => x"dcce7b00",
   400 => x"18183000",
   401 => x"00000000",
   402 => x"0c183030",
   403 => x"30180c00",
   404 => x"30180c0c",
   405 => x"0c183000",
   406 => x"00663cff",
   407 => x"3c660000",
   408 => x"0018187e",
   409 => x"18180000",
   410 => x"00000000",
   411 => x"00181830",
   412 => x"0000007e",
   413 => x"00000000",
   414 => x"00000000",
   415 => x"00181800",
   416 => x"03060c18",
   417 => x"3060c000",
   418 => x"3c666e7e",
   419 => x"76663c00",
   420 => x"18387818",
   421 => x"18181800",
   422 => x"3c66060c",
   423 => x"18307e00",
   424 => x"3c66061c",
   425 => x"06663c00",
   426 => x"1c3c6ccc",
   427 => x"fe0c0c00",
   428 => x"7e607c06",
   429 => x"06663c00",
   430 => x"1c30607c",
   431 => x"66663c00",
   432 => x"7e06060c",
   433 => x"18181800",
   434 => x"3c66663c",
   435 => x"66663c00",
   436 => x"3c66663e",
   437 => x"060c3800",
   438 => x"00181800",
   439 => x"00181800",
   440 => x"00181800",
   441 => x"00181830",
   442 => x"00061860",
   443 => x"18060000",
   444 => x"00007e00",
   445 => x"7e000000",
   446 => x"00601806",
   447 => x"18600000",
   448 => x"3c66060c",
   449 => x"18001800",
   450 => x"7cc6ded6",
   451 => x"dec07800",
   452 => x"3c66667e",
   453 => x"66666600",
   454 => x"7c66667c",
   455 => x"66667c00",
   456 => x"1e306060",
   457 => x"60301e00",
   458 => x"786c6666",
   459 => x"666c7800",
   460 => x"7e606078",
   461 => x"60607e00",
   462 => x"7e606078",
   463 => x"60606000",
   464 => x"3c66606e",
   465 => x"66663e00",
   466 => x"6666667e",
   467 => x"66666600",
   468 => x"3c181818",
   469 => x"18183c00",
   470 => x"06060606",
   471 => x"06663c00",
   472 => x"c6ccd8f0",
   473 => x"d8ccc600",
   474 => x"60606060",
   475 => x"60607e00",
   476 => x"c6eefed6",
   477 => x"c6c6c600",
   478 => x"c6e6f6de",
   479 => x"cec6c600",
   480 => x"3c666666",
   481 => x"66663c00",
   482 => x"7c66667c",
   483 => x"60606000",
   484 => x"78cccccc",
   485 => x"ccdc7e00",
   486 => x"7c66667c",
   487 => x"6c666600",
   488 => x"3c66703c",
   489 => x"0e663c00",
   490 => x"7e181818",
   491 => x"18181800",
   492 => x"66666666",
   493 => x"66663c00",
   494 => x"66666666",
   495 => x"3c3c1800",
   496 => x"c6c6c6d6",
   497 => x"feeec600",
   498 => x"c3663c18",
   499 => x"3c66c300",
   500 => x"c3663c18",
   501 => x"18181800",
   502 => x"fe0c1830",
   503 => x"60c0fe00",
   504 => x"3c303030",
   505 => x"30303c00",
   506 => x"c0603018",
   507 => x"0c060300",
   508 => x"3c0c0c0c",
   509 => x"0c0c3c00",
   510 => x"10386cc6",
   511 => x"00000000",
   512 => x"00000000",
   513 => x"000000fe",
   514 => x"18180c00",
   515 => x"00000000",
   516 => x"00003c06",
   517 => x"3e663e00",
   518 => x"60607c66",
   519 => x"66667c00",
   520 => x"00003c60",
   521 => x"60603c00",
   522 => x"06063e66",
   523 => x"66663e00",
   524 => x"00003c66",
   525 => x"7e603c00",
   526 => x"1c307c30",
   527 => x"30303000",
   528 => x"00003e66",
   529 => x"663e063c",
   530 => x"60607c66",
   531 => x"66666600",
   532 => x"18001818",
   533 => x"18180c00",
   534 => x"0c000c0c",
   535 => x"0c0c0c78",
   536 => x"6060666c",
   537 => x"786c6600",
   538 => x"18181818",
   539 => x"18180c00",
   540 => x"0000ecfe",
   541 => x"d6c6c600",
   542 => x"00007c66",
   543 => x"66666600",
   544 => x"00003c66",
   545 => x"66663c00",
   546 => x"00007c66",
   547 => x"667c6060",
   548 => x"00003e66",
   549 => x"663e0606",
   550 => x"00007c66",
   551 => x"60606000",
   552 => x"00003c60",
   553 => x"3c067c00",
   554 => x"30307c30",
   555 => x"30301c00",
   556 => x"00006666",
   557 => x"66663e00",
   558 => x"00006666",
   559 => x"663c1800",
   560 => x"0000c6c6",
   561 => x"d6fe6c00",
   562 => x"0000c66c",
   563 => x"386cc600",
   564 => x"00006666",
   565 => x"663c1830",
   566 => x"00007e0c",
   567 => x"18307e00",
   568 => x"0e181870",
   569 => x"18180e00",
   570 => x"18181818",
   571 => x"18181800",
   572 => x"7018180e",
   573 => x"18187000",
   574 => x"729c0000",
   575 => x"00000000",
   576 => x"fefefefe",
   577 => x"fefefe00",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
   785 => x"00000000",
   786 => x"00000000",
   787 => x"00000000",
   788 => x"00000000",
   789 => x"00000000",
   790 => x"00000000",
   791 => x"00000000",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
   799 => x"00000000",
   800 => x"00000000",
   801 => x"00000000",
   802 => x"00000000",
   803 => x"00000000",
   804 => x"00000000",
   805 => x"00000000",
   806 => x"00000000",
   807 => x"00000000",
   808 => x"00000000",
   809 => x"00000000",
   810 => x"00000000",
   811 => x"00000000",
   812 => x"00000000",
   813 => x"00000000",
   814 => x"00000000",
   815 => x"00000000",
   816 => x"00000000",
   817 => x"00000000",
   818 => x"00000000",
   819 => x"00000000",
   820 => x"00000000",
   821 => x"00000000",
   822 => x"00000000",
   823 => x"00000000",
   824 => x"00000000",
   825 => x"00000000",
   826 => x"00000000",
   827 => x"00000000",
   828 => x"00000000",
   829 => x"00000000",
   830 => x"00000000",
   831 => x"00000000",
   832 => x"00000000",
   833 => x"00000000",
   834 => x"30313233",
   835 => x"34353637",
   836 => x"38394142",
   837 => x"43444546",
   838 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

