-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"80700b0b",
     2 => x"80c9a80c",
     3 => x"3a0b0b0b",
     4 => x"b9e20400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"8f040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80c4",
   162 => x"d0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f7040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"df040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80c9a40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"83e23fbc",
   257 => x"9e3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104b0",
   280 => x"08b408b8",
   281 => x"0875759e",
   282 => x"f62d5050",
   283 => x"b00856b8",
   284 => x"0cb40cb0",
   285 => x"0c5104b0",
   286 => x"08b408b8",
   287 => x"0875759d",
   288 => x"c42d5050",
   289 => x"b00856b8",
   290 => x"0cb40cb0",
   291 => x"0c5104b0",
   292 => x"08b408b8",
   293 => x"08baa92d",
   294 => x"b80cb40c",
   295 => x"b00c04fe",
   296 => x"3d0d0b0b",
   297 => x"80e79408",
   298 => x"53841308",
   299 => x"70882a70",
   300 => x"81065152",
   301 => x"5270802e",
   302 => x"f0387181",
   303 => x"ff06b00c",
   304 => x"843d0d04",
   305 => x"ff3d0d0b",
   306 => x"0b80e794",
   307 => x"08527108",
   308 => x"70882a81",
   309 => x"32708106",
   310 => x"51515170",
   311 => x"f1387372",
   312 => x"0c833d0d",
   313 => x"0480c9a4",
   314 => x"08802ea4",
   315 => x"3880c9a8",
   316 => x"08822ebd",
   317 => x"38838080",
   318 => x"0b0b0b80",
   319 => x"e7940c82",
   320 => x"a0800b80",
   321 => x"e7980c82",
   322 => x"90800b80",
   323 => x"e79c0c04",
   324 => x"f8808080",
   325 => x"a40b0b0b",
   326 => x"80e7940c",
   327 => x"f8808082",
   328 => x"800b80e7",
   329 => x"980cf880",
   330 => x"8084800b",
   331 => x"80e79c0c",
   332 => x"0480c0a8",
   333 => x"808c0b0b",
   334 => x"0b80e794",
   335 => x"0c80c0a8",
   336 => x"80940b80",
   337 => x"e7980c80",
   338 => x"c4e00b80",
   339 => x"e79c0c04",
   340 => x"f23d0d60",
   341 => x"80e79808",
   342 => x"565d8275",
   343 => x"0c805980",
   344 => x"5a800b8f",
   345 => x"3d5d5b7a",
   346 => x"10101570",
   347 => x"08710871",
   348 => x"9f2c7e85",
   349 => x"2b585555",
   350 => x"7d535957",
   351 => x"90d03f7d",
   352 => x"7f7a7207",
   353 => x"7c720771",
   354 => x"71608105",
   355 => x"415f5d5b",
   356 => x"59575581",
   357 => x"7b278f38",
   358 => x"767d0c77",
   359 => x"841e0c7c",
   360 => x"b00c903d",
   361 => x"0d0480e7",
   362 => x"980855ff",
   363 => x"ba39ff3d",
   364 => x"0d80e7a0",
   365 => x"335170a7",
   366 => x"3880c9b0",
   367 => x"08700852",
   368 => x"5270802e",
   369 => x"94388412",
   370 => x"80c9b00c",
   371 => x"702d80c9",
   372 => x"b0087008",
   373 => x"525270ee",
   374 => x"38810b80",
   375 => x"e7a03483",
   376 => x"3d0d0404",
   377 => x"803d0d0b",
   378 => x"0b80e790",
   379 => x"08802e8e",
   380 => x"380b0b0b",
   381 => x"0b800b80",
   382 => x"2e098106",
   383 => x"8538823d",
   384 => x"0d040b0b",
   385 => x"80e79051",
   386 => x"0b0b0bf3",
   387 => x"f33f823d",
   388 => x"0d0404f7",
   389 => x"3d0d7c84",
   390 => x"11085555",
   391 => x"817c25b9",
   392 => x"387351a3",
   393 => x"e33f873d",
   394 => x"7054b008",
   395 => x"53745256",
   396 => x"81883f80",
   397 => x"55741670",
   398 => x"33535480",
   399 => x"c4f8518c",
   400 => x"983f8115",
   401 => x"558f7525",
   402 => x"ec3880c9",
   403 => x"90518b99",
   404 => x"3f800bb0",
   405 => x"0c8b3d0d",
   406 => x"04740852",
   407 => x"80c4e451",
   408 => x"8bf73f81",
   409 => x"0bb00c8b",
   410 => x"3d0d04fe",
   411 => x"3d0d7476",
   412 => x"54527173",
   413 => x"3471882a",
   414 => x"51708114",
   415 => x"3471902a",
   416 => x"51708214",
   417 => x"3471982a",
   418 => x"52718314",
   419 => x"34843d0d",
   420 => x"04fd3d0d",
   421 => x"75811133",
   422 => x"71337188",
   423 => x"2b078213",
   424 => x"3370902b",
   425 => x"72078315",
   426 => x"3370982b",
   427 => x"7207b00c",
   428 => x"55525253",
   429 => x"5452853d",
   430 => x"0d04da3d",
   431 => x"0daa3d08",
   432 => x"ac3d0848",
   433 => x"5786ba94",
   434 => x"c68143fe",
   435 => x"feb6d789",
   436 => x"44f9c5eb",
   437 => x"b9fe4581",
   438 => x"81c9a8f6",
   439 => x"0b811870",
   440 => x"71bf0657",
   441 => x"57414673",
   442 => x"b82e9138",
   443 => x"7f810570",
   444 => x"bf065540",
   445 => x"73b82e09",
   446 => x"8106f138",
   447 => x"7f880551",
   448 => x"94a03fb0",
   449 => x"087754aa",
   450 => x"3d0853b0",
   451 => x"085242a0",
   452 => x"a83f6117",
   453 => x"56ff8076",
   454 => x"34746027",
   455 => x"8f386115",
   456 => x"58807834",
   457 => x"8115557f",
   458 => x"7526f338",
   459 => x"76832b62",
   460 => x"61055a5b",
   461 => x"7a79347a",
   462 => x"882a5d7c",
   463 => x"811a347a",
   464 => x"902a5c7b",
   465 => x"821a347a",
   466 => x"982a5a79",
   467 => x"831a3476",
   468 => x"9d2a841a",
   469 => x"58557477",
   470 => x"34800b81",
   471 => x"1834800b",
   472 => x"82183480",
   473 => x"0b831834",
   474 => x"80416060",
   475 => x"2781be38",
   476 => x"800b993d",
   477 => x"63630557",
   478 => x"58568115",
   479 => x"33753371",
   480 => x"882b0782",
   481 => x"17337090",
   482 => x"2b720783",
   483 => x"19337098",
   484 => x"2b72077c",
   485 => x"7084055e",
   486 => x"0c434181",
   487 => x"19841959",
   488 => x"595a555a",
   489 => x"8f7627d2",
   490 => x"38626466",
   491 => x"685d5a56",
   492 => x"5f80705f",
   493 => x"59855d81",
   494 => x"5c788f26",
   495 => x"81f93874",
   496 => x"097a0675",
   497 => x"79060779",
   498 => x"57577882",
   499 => x"2b547978",
   500 => x"76611a80",
   501 => x"c7801808",
   502 => x"05ac3d7a",
   503 => x"10100580",
   504 => x"c5801908",
   505 => x"c0120813",
   506 => x"c0130814",
   507 => x"a073312a",
   508 => x"71732b07",
   509 => x"75057761",
   510 => x"81056585",
   511 => x"05678305",
   512 => x"6987054a",
   513 => x"48464247",
   514 => x"545a5c5a",
   515 => x"585a5b5b",
   516 => x"bf7927ff",
   517 => x"a438621b",
   518 => x"6416661a",
   519 => x"681d6480",
   520 => x"c0054549",
   521 => x"4745437f",
   522 => x"6126fec4",
   523 => x"38615192",
   524 => x"813f6267",
   525 => x"3462882a",
   526 => x"55746781",
   527 => x"05346290",
   528 => x"2a577667",
   529 => x"82053462",
   530 => x"982a5473",
   531 => x"67830534",
   532 => x"66840558",
   533 => x"63783463",
   534 => x"882a5b7a",
   535 => x"81193463",
   536 => x"902a5a79",
   537 => x"82193463",
   538 => x"982a5978",
   539 => x"83193466",
   540 => x"88054464",
   541 => x"64346488",
   542 => x"2a5e7d64",
   543 => x"81053464",
   544 => x"902a5d7c",
   545 => x"64820534",
   546 => x"64982a5c",
   547 => x"7b648305",
   548 => x"34668c05",
   549 => x"40656034",
   550 => x"65882a43",
   551 => x"62608105",
   552 => x"3465902a",
   553 => x"42616082",
   554 => x"05346598",
   555 => x"2a416060",
   556 => x"830534a8",
   557 => x"3d0d0478",
   558 => x"9f2680db",
   559 => x"38790978",
   560 => x"067a7606",
   561 => x"0779822b",
   562 => x"7d8f067c",
   563 => x"7b795d5e",
   564 => x"5e58557f",
   565 => x"0580c780",
   566 => x"150805a9",
   567 => x"3d771010",
   568 => x"0580c580",
   569 => x"1608c012",
   570 => x"0813c013",
   571 => x"0814a073",
   572 => x"312a7173",
   573 => x"2b077c05",
   574 => x"7f811f62",
   575 => x"85056483",
   576 => x"05668705",
   577 => x"4745435f",
   578 => x"44545759",
   579 => x"5755bf79",
   580 => x"27fda638",
   581 => x"fe803974",
   582 => x"78327a32",
   583 => x"7d8f0657",
   584 => x"57af7927",
   585 => x"fda43879",
   586 => x"09750778",
   587 => x"327e8f06",
   588 => x"7a822b56",
   589 => x"5757fd96",
   590 => x"39ff3d0d",
   591 => x"fea0800b",
   592 => x"86ffe280",
   593 => x"23800b86",
   594 => x"ffe28223",
   595 => x"800b86ff",
   596 => x"e2842380",
   597 => x"0b86ffe2",
   598 => x"8823800b",
   599 => x"86ffe28a",
   600 => x"23828080",
   601 => x"52a0bf51",
   602 => x"80727084",
   603 => x"05540cff",
   604 => x"11517080",
   605 => x"25f238bc",
   606 => x"0b86ffe1",
   607 => x"922381d4",
   608 => x"0b86ffe1",
   609 => x"942380d9",
   610 => x"810b86ff",
   611 => x"e18e23e9",
   612 => x"c10b86ff",
   613 => x"e1902386",
   614 => x"ff0b86ff",
   615 => x"e380239f",
   616 => x"ff0b86ff",
   617 => x"e3822380",
   618 => x"d7b40870",
   619 => x"535181e0",
   620 => x"72708205",
   621 => x"54238072",
   622 => x"70820554",
   623 => x"2381e272",
   624 => x"70820554",
   625 => x"23fe8080",
   626 => x"72708205",
   627 => x"5423ff72",
   628 => x"70820554",
   629 => x"23fe7223",
   630 => x"70902c52",
   631 => x"7186ffe1",
   632 => x"80237086",
   633 => x"ffe18223",
   634 => x"800b86ff",
   635 => x"e18823fe",
   636 => x"87900b86",
   637 => x"ffe19623",
   638 => x"800b80e7",
   639 => x"a40c800b",
   640 => x"80e7a80c",
   641 => x"833d0d04",
   642 => x"fb3d0d02",
   643 => x"9f053380",
   644 => x"e7a808b1",
   645 => x"800a2980",
   646 => x"e7a40805",
   647 => x"71a02916",
   648 => x"f8801108",
   649 => x"f8841208",
   650 => x"52575754",
   651 => x"56737334",
   652 => x"73ffb014",
   653 => x"3473fee0",
   654 => x"143473fe",
   655 => x"90143474",
   656 => x"fdc01434",
   657 => x"74fcf014",
   658 => x"3474fca0",
   659 => x"143474fb",
   660 => x"d0143475",
   661 => x"8a2e80e8",
   662 => x"3880e7a4",
   663 => x"08810580",
   664 => x"e7a40c80",
   665 => x"e7a40880",
   666 => x"d02eb638",
   667 => x"80e7a808",
   668 => x"992e8538",
   669 => x"873d0d04",
   670 => x"82808055",
   671 => x"82858054",
   672 => x"9f9f5373",
   673 => x"70840555",
   674 => x"08757084",
   675 => x"05570cff",
   676 => x"13537280",
   677 => x"25ed3898",
   678 => x"0b80e7a8",
   679 => x"0c873d0d",
   680 => x"0480e7a8",
   681 => x"08810580",
   682 => x"e7a80c80",
   683 => x"0b80e7a4",
   684 => x"0c80e7a8",
   685 => x"08992e09",
   686 => x"8106ffb8",
   687 => x"38ffb939",
   688 => x"80e7a808",
   689 => x"810580e7",
   690 => x"a80c80e7",
   691 => x"a808992e",
   692 => x"098106ff",
   693 => x"9f38ffa0",
   694 => x"39f83d0d",
   695 => x"7a707081",
   696 => x"05523358",
   697 => x"5976802e",
   698 => x"80f43880",
   699 => x"e7a808b1",
   700 => x"800a2980",
   701 => x"e7a40805",
   702 => x"77a02919",
   703 => x"f8801108",
   704 => x"f8841208",
   705 => x"5957f888",
   706 => x"05595474",
   707 => x"743474ff",
   708 => x"b0153474",
   709 => x"fee01534",
   710 => x"74fe9015",
   711 => x"3475fdc0",
   712 => x"153475fc",
   713 => x"f0153475",
   714 => x"fca01534",
   715 => x"75fbd015",
   716 => x"34768a2e",
   717 => x"80f93880",
   718 => x"e7a40881",
   719 => x"0580e7a4",
   720 => x"0c80e7a4",
   721 => x"0880d02e",
   722 => x"80c63880",
   723 => x"e7a80899",
   724 => x"2e903878",
   725 => x"7081055a",
   726 => x"335776ff",
   727 => x"8e388a3d",
   728 => x"0d048280",
   729 => x"80558285",
   730 => x"80549f9f",
   731 => x"53737084",
   732 => x"05550875",
   733 => x"70840557",
   734 => x"0cff1353",
   735 => x"728025ed",
   736 => x"38980b80",
   737 => x"e7a80c78",
   738 => x"7081055a",
   739 => x"3357cb39",
   740 => x"80e7a808",
   741 => x"810580e7",
   742 => x"a80c800b",
   743 => x"80e7a40c",
   744 => x"80e7a808",
   745 => x"992e0981",
   746 => x"06ffa838",
   747 => x"ffb43980",
   748 => x"e7a80881",
   749 => x"0580e7a8",
   750 => x"0c80e7a8",
   751 => x"08992e09",
   752 => x"8106ff8f",
   753 => x"38ff9b39",
   754 => x"ff3d0d02",
   755 => x"8f053352",
   756 => x"ff840870",
   757 => x"882a7081",
   758 => x"06515151",
   759 => x"70802ef0",
   760 => x"3871ff84",
   761 => x"0c833d0d",
   762 => x"04fe3d0d",
   763 => x"74703352",
   764 => x"5370802e",
   765 => x"a1387052",
   766 => x"811353ff",
   767 => x"84087088",
   768 => x"2a708106",
   769 => x"51515170",
   770 => x"802ef038",
   771 => x"71ff840c",
   772 => x"72335271",
   773 => x"e338843d",
   774 => x"0d04ff3d",
   775 => x"0dff8408",
   776 => x"70892a70",
   777 => x"81065152",
   778 => x"5270802e",
   779 => x"f0387181",
   780 => x"ff06b00c",
   781 => x"833d0d04",
   782 => x"ff3d0d02",
   783 => x"8f053352",
   784 => x"ff840870",
   785 => x"882a7081",
   786 => x"06515151",
   787 => x"70802ef0",
   788 => x"3871ff84",
   789 => x"0c833d0d",
   790 => x"04f53d0d",
   791 => x"8e3d7070",
   792 => x"84055208",
   793 => x"98b85b55",
   794 => x"5b807470",
   795 => x"81055633",
   796 => x"755a5457",
   797 => x"72772ebe",
   798 => x"3872a52e",
   799 => x"09810680",
   800 => x"c5387770",
   801 => x"81055933",
   802 => x"537280e4",
   803 => x"2e81b638",
   804 => x"7280e424",
   805 => x"80c63872",
   806 => x"80e32ea1",
   807 => x"388052a5",
   808 => x"51782d80",
   809 => x"52725178",
   810 => x"2d821757",
   811 => x"77708105",
   812 => x"59335372",
   813 => x"c43876b0",
   814 => x"0c8d3d0d",
   815 => x"047a841c",
   816 => x"83123355",
   817 => x"5c568052",
   818 => x"7251782d",
   819 => x"81177870",
   820 => x"81055a33",
   821 => x"545772ff",
   822 => x"a038db39",
   823 => x"7280f32e",
   824 => x"098106ff",
   825 => x"b8387a84",
   826 => x"1c710858",
   827 => x"5c548076",
   828 => x"335b5579",
   829 => x"752e8d38",
   830 => x"81157017",
   831 => x"7033555b",
   832 => x"5572f538",
   833 => x"ff155480",
   834 => x"7525ffa0",
   835 => x"38757081",
   836 => x"05573353",
   837 => x"80527251",
   838 => x"782d8117",
   839 => x"74ff1656",
   840 => x"56578075",
   841 => x"25ff8538",
   842 => x"75708105",
   843 => x"57335380",
   844 => x"52725178",
   845 => x"2d811774",
   846 => x"ff165656",
   847 => x"57748024",
   848 => x"cc38fee8",
   849 => x"397a841c",
   850 => x"710880e8",
   851 => x"840b80e7",
   852 => x"ac545d56",
   853 => x"5c558056",
   854 => x"73762e09",
   855 => x"8106b838",
   856 => x"b00b80e7",
   857 => x"ac348115",
   858 => x"55ff1555",
   859 => x"74337a70",
   860 => x"81055c34",
   861 => x"81165674",
   862 => x"80e7ac2e",
   863 => x"098106e9",
   864 => x"38807a34",
   865 => x"7580e884",
   866 => x"0bff1256",
   867 => x"57557480",
   868 => x"24fefa38",
   869 => x"fe963973",
   870 => x"8f0680c9",
   871 => x"80055372",
   872 => x"33757081",
   873 => x"05573473",
   874 => x"842a5473",
   875 => x"ea387480",
   876 => x"e7ac2ecd",
   877 => x"38ff1555",
   878 => x"74337a70",
   879 => x"81055c34",
   880 => x"81165674",
   881 => x"80e7ac2e",
   882 => x"ffb738ff",
   883 => x"9c39bc08",
   884 => x"02bc0cf5",
   885 => x"3d0dbc08",
   886 => x"9405089d",
   887 => x"38bc088c",
   888 => x"0508bc08",
   889 => x"900508bc",
   890 => x"08880508",
   891 => x"58565473",
   892 => x"760c7484",
   893 => x"170c81bf",
   894 => x"39800bbc",
   895 => x"08f0050c",
   896 => x"800bbc08",
   897 => x"f4050cbc",
   898 => x"088c0508",
   899 => x"bc089005",
   900 => x"08565473",
   901 => x"bc08f005",
   902 => x"0c74bc08",
   903 => x"f4050cbc",
   904 => x"08f805bc",
   905 => x"08f00556",
   906 => x"56887054",
   907 => x"75537652",
   908 => x"5492863f",
   909 => x"a00bbc08",
   910 => x"94050831",
   911 => x"bc08ec05",
   912 => x"0cbc08ec",
   913 => x"05088024",
   914 => x"9d38800b",
   915 => x"bc08f405",
   916 => x"0cbc08ec",
   917 => x"050830bc",
   918 => x"08fc0508",
   919 => x"712bbc08",
   920 => x"f0050c54",
   921 => x"b939bc08",
   922 => x"fc0508bc",
   923 => x"08ec0508",
   924 => x"2abc08e8",
   925 => x"050cbc08",
   926 => x"fc0508bc",
   927 => x"08940508",
   928 => x"2bbc08f4",
   929 => x"050cbc08",
   930 => x"f80508bc",
   931 => x"08940508",
   932 => x"2b70bc08",
   933 => x"e8050807",
   934 => x"bc08f005",
   935 => x"0c54bc08",
   936 => x"f00508bc",
   937 => x"08f40508",
   938 => x"bc088805",
   939 => x"08585654",
   940 => x"73760c74",
   941 => x"84170cbc",
   942 => x"08880508",
   943 => x"b00c8d3d",
   944 => x"0dbc0c04",
   945 => x"bc0802bc",
   946 => x"0cf93d0d",
   947 => x"800bbc08",
   948 => x"fc050cbc",
   949 => x"08880508",
   950 => x"8025ab38",
   951 => x"bc088805",
   952 => x"0830bc08",
   953 => x"88050c80",
   954 => x"0bbc08f4",
   955 => x"050cbc08",
   956 => x"fc050888",
   957 => x"38810bbc",
   958 => x"08f4050c",
   959 => x"bc08f405",
   960 => x"08bc08fc",
   961 => x"050cbc08",
   962 => x"8c050880",
   963 => x"25ab38bc",
   964 => x"088c0508",
   965 => x"30bc088c",
   966 => x"050c800b",
   967 => x"bc08f005",
   968 => x"0cbc08fc",
   969 => x"05088838",
   970 => x"810bbc08",
   971 => x"f0050cbc",
   972 => x"08f00508",
   973 => x"bc08fc05",
   974 => x"0c8053bc",
   975 => x"088c0508",
   976 => x"52bc0888",
   977 => x"05085181",
   978 => x"a73fb008",
   979 => x"70bc08f8",
   980 => x"050c54bc",
   981 => x"08fc0508",
   982 => x"802e8c38",
   983 => x"bc08f805",
   984 => x"0830bc08",
   985 => x"f8050cbc",
   986 => x"08f80508",
   987 => x"70b00c54",
   988 => x"893d0dbc",
   989 => x"0c04bc08",
   990 => x"02bc0cfb",
   991 => x"3d0d800b",
   992 => x"bc08fc05",
   993 => x"0cbc0888",
   994 => x"05088025",
   995 => x"9338bc08",
   996 => x"88050830",
   997 => x"bc088805",
   998 => x"0c810bbc",
   999 => x"08fc050c",
  1000 => x"bc088c05",
  1001 => x"0880258c",
  1002 => x"38bc088c",
  1003 => x"050830bc",
  1004 => x"088c050c",
  1005 => x"8153bc08",
  1006 => x"8c050852",
  1007 => x"bc088805",
  1008 => x"0851ad3f",
  1009 => x"b00870bc",
  1010 => x"08f8050c",
  1011 => x"54bc08fc",
  1012 => x"0508802e",
  1013 => x"8c38bc08",
  1014 => x"f8050830",
  1015 => x"bc08f805",
  1016 => x"0cbc08f8",
  1017 => x"050870b0",
  1018 => x"0c54873d",
  1019 => x"0dbc0c04",
  1020 => x"bc0802bc",
  1021 => x"0cfd3d0d",
  1022 => x"810bbc08",
  1023 => x"fc050c80",
  1024 => x"0bbc08f8",
  1025 => x"050cbc08",
  1026 => x"8c0508bc",
  1027 => x"08880508",
  1028 => x"27ac38bc",
  1029 => x"08fc0508",
  1030 => x"802ea338",
  1031 => x"800bbc08",
  1032 => x"8c050824",
  1033 => x"9938bc08",
  1034 => x"8c050810",
  1035 => x"bc088c05",
  1036 => x"0cbc08fc",
  1037 => x"050810bc",
  1038 => x"08fc050c",
  1039 => x"c939bc08",
  1040 => x"fc050880",
  1041 => x"2e80c938",
  1042 => x"bc088c05",
  1043 => x"08bc0888",
  1044 => x"050826a1",
  1045 => x"38bc0888",
  1046 => x"0508bc08",
  1047 => x"8c050831",
  1048 => x"bc088805",
  1049 => x"0cbc08f8",
  1050 => x"0508bc08",
  1051 => x"fc050807",
  1052 => x"bc08f805",
  1053 => x"0cbc08fc",
  1054 => x"0508812a",
  1055 => x"bc08fc05",
  1056 => x"0cbc088c",
  1057 => x"0508812a",
  1058 => x"bc088c05",
  1059 => x"0cffaf39",
  1060 => x"bc089005",
  1061 => x"08802e8f",
  1062 => x"38bc0888",
  1063 => x"050870bc",
  1064 => x"08f4050c",
  1065 => x"518d39bc",
  1066 => x"08f80508",
  1067 => x"70bc08f4",
  1068 => x"050c51bc",
  1069 => x"08f40508",
  1070 => x"b00c853d",
  1071 => x"0dbc0c04",
  1072 => x"bc0802bc",
  1073 => x"0cff3d0d",
  1074 => x"800bbc08",
  1075 => x"fc050cbc",
  1076 => x"08880508",
  1077 => x"8106ff11",
  1078 => x"700970bc",
  1079 => x"088c0508",
  1080 => x"06bc08fc",
  1081 => x"050811bc",
  1082 => x"08fc050c",
  1083 => x"bc088805",
  1084 => x"08812abc",
  1085 => x"0888050c",
  1086 => x"bc088c05",
  1087 => x"0810bc08",
  1088 => x"8c050c51",
  1089 => x"515151bc",
  1090 => x"08880508",
  1091 => x"802e8438",
  1092 => x"ffbd39bc",
  1093 => x"08fc0508",
  1094 => x"70b00c51",
  1095 => x"833d0dbc",
  1096 => x"0c04ff3d",
  1097 => x"0d735280",
  1098 => x"dffc0851",
  1099 => x"963f833d",
  1100 => x"0d04ff3d",
  1101 => x"0d735280",
  1102 => x"dffc0851",
  1103 => x"8fdf3f83",
  1104 => x"3d0d04f3",
  1105 => x"3d0d7f61",
  1106 => x"8b1170f8",
  1107 => x"065c5555",
  1108 => x"5e729626",
  1109 => x"83389059",
  1110 => x"80792474",
  1111 => x"7a260753",
  1112 => x"80547274",
  1113 => x"2e098106",
  1114 => x"80cb387d",
  1115 => x"518ce33f",
  1116 => x"7883f726",
  1117 => x"80c63878",
  1118 => x"832a7010",
  1119 => x"101080d7",
  1120 => x"f4058c11",
  1121 => x"0859595a",
  1122 => x"76782e83",
  1123 => x"b0388417",
  1124 => x"08fc0656",
  1125 => x"8c170888",
  1126 => x"1808718c",
  1127 => x"120c8812",
  1128 => x"0c587517",
  1129 => x"84110881",
  1130 => x"0784120c",
  1131 => x"537d518c",
  1132 => x"a23f8817",
  1133 => x"5473b00c",
  1134 => x"8f3d0d04",
  1135 => x"78892a79",
  1136 => x"832a5b53",
  1137 => x"72802ebf",
  1138 => x"3878862a",
  1139 => x"b8055a84",
  1140 => x"7327b438",
  1141 => x"80db135a",
  1142 => x"947327ab",
  1143 => x"38788c2a",
  1144 => x"80ee055a",
  1145 => x"80d47327",
  1146 => x"9e38788f",
  1147 => x"2a80f705",
  1148 => x"5a82d473",
  1149 => x"27913878",
  1150 => x"922a80fc",
  1151 => x"055a8ad4",
  1152 => x"73278438",
  1153 => x"80fe5a79",
  1154 => x"10101080",
  1155 => x"d7f4058c",
  1156 => x"11085855",
  1157 => x"76752ea3",
  1158 => x"38841708",
  1159 => x"fc06707a",
  1160 => x"31555673",
  1161 => x"8f2488d5",
  1162 => x"38738025",
  1163 => x"fee6388c",
  1164 => x"17085776",
  1165 => x"752e0981",
  1166 => x"06df3881",
  1167 => x"1a5a80d8",
  1168 => x"84085776",
  1169 => x"80d7fc2e",
  1170 => x"82c03884",
  1171 => x"1708fc06",
  1172 => x"707a3155",
  1173 => x"56738f24",
  1174 => x"81f93880",
  1175 => x"d7fc0b80",
  1176 => x"d8880c80",
  1177 => x"d7fc0b80",
  1178 => x"d8840c73",
  1179 => x"8025feb2",
  1180 => x"3883ff76",
  1181 => x"2783df38",
  1182 => x"75892a76",
  1183 => x"832a5553",
  1184 => x"72802ebf",
  1185 => x"3875862a",
  1186 => x"b8055484",
  1187 => x"7327b438",
  1188 => x"80db1354",
  1189 => x"947327ab",
  1190 => x"38758c2a",
  1191 => x"80ee0554",
  1192 => x"80d47327",
  1193 => x"9e38758f",
  1194 => x"2a80f705",
  1195 => x"5482d473",
  1196 => x"27913875",
  1197 => x"922a80fc",
  1198 => x"05548ad4",
  1199 => x"73278438",
  1200 => x"80fe5473",
  1201 => x"10101080",
  1202 => x"d7f40588",
  1203 => x"11085658",
  1204 => x"74782e86",
  1205 => x"cf388415",
  1206 => x"08fc0653",
  1207 => x"7573278d",
  1208 => x"38881508",
  1209 => x"5574782e",
  1210 => x"098106ea",
  1211 => x"388c1508",
  1212 => x"80d7f40b",
  1213 => x"84050871",
  1214 => x"8c1a0c76",
  1215 => x"881a0c78",
  1216 => x"88130c78",
  1217 => x"8c180c5d",
  1218 => x"58795380",
  1219 => x"7a2483e6",
  1220 => x"3872822c",
  1221 => x"81712b5c",
  1222 => x"537a7c26",
  1223 => x"8198387b",
  1224 => x"7b065372",
  1225 => x"82f13879",
  1226 => x"fc068405",
  1227 => x"5a7a1070",
  1228 => x"7d06545b",
  1229 => x"7282e038",
  1230 => x"841a5af1",
  1231 => x"3988178c",
  1232 => x"11085858",
  1233 => x"76782e09",
  1234 => x"8106fcc2",
  1235 => x"38821a5a",
  1236 => x"fdec3978",
  1237 => x"17798107",
  1238 => x"84190c70",
  1239 => x"80d8880c",
  1240 => x"7080d884",
  1241 => x"0c80d7fc",
  1242 => x"0b8c120c",
  1243 => x"8c110888",
  1244 => x"120c7481",
  1245 => x"0784120c",
  1246 => x"74117571",
  1247 => x"0c51537d",
  1248 => x"5188d03f",
  1249 => x"881754fc",
  1250 => x"ac3980d7",
  1251 => x"f40b8405",
  1252 => x"087a545c",
  1253 => x"798025fe",
  1254 => x"f83882da",
  1255 => x"397a097c",
  1256 => x"067080d7",
  1257 => x"f40b8405",
  1258 => x"0c5c7a10",
  1259 => x"5b7a7c26",
  1260 => x"85387a85",
  1261 => x"b83880d7",
  1262 => x"f40b8805",
  1263 => x"08708412",
  1264 => x"08fc0670",
  1265 => x"7c317c72",
  1266 => x"268f7225",
  1267 => x"0757575c",
  1268 => x"5d557280",
  1269 => x"2e80db38",
  1270 => x"797a1680",
  1271 => x"d7ec081b",
  1272 => x"90115a55",
  1273 => x"575b80d7",
  1274 => x"e808ff2e",
  1275 => x"8838a08f",
  1276 => x"13e08006",
  1277 => x"5776527d",
  1278 => x"5187d93f",
  1279 => x"b00854b0",
  1280 => x"08ff2e90",
  1281 => x"38b00876",
  1282 => x"27829938",
  1283 => x"7480d7f4",
  1284 => x"2e829138",
  1285 => x"80d7f40b",
  1286 => x"88050855",
  1287 => x"841508fc",
  1288 => x"06707a31",
  1289 => x"7a72268f",
  1290 => x"72250752",
  1291 => x"55537283",
  1292 => x"e6387479",
  1293 => x"81078417",
  1294 => x"0c791670",
  1295 => x"80d7f40b",
  1296 => x"88050c75",
  1297 => x"81078412",
  1298 => x"0c547e52",
  1299 => x"5787843f",
  1300 => x"881754fa",
  1301 => x"e0397583",
  1302 => x"2a705454",
  1303 => x"80742481",
  1304 => x"9b387282",
  1305 => x"2c81712b",
  1306 => x"80d7f808",
  1307 => x"077080d7",
  1308 => x"f40b8405",
  1309 => x"0c751010",
  1310 => x"1080d7f4",
  1311 => x"05881108",
  1312 => x"585a5d53",
  1313 => x"778c180c",
  1314 => x"7488180c",
  1315 => x"7688190c",
  1316 => x"768c160c",
  1317 => x"fcf33979",
  1318 => x"7a101010",
  1319 => x"80d7f405",
  1320 => x"7057595d",
  1321 => x"8c150857",
  1322 => x"76752ea3",
  1323 => x"38841708",
  1324 => x"fc06707a",
  1325 => x"31555673",
  1326 => x"8f2483ca",
  1327 => x"38738025",
  1328 => x"8481388c",
  1329 => x"17085776",
  1330 => x"752e0981",
  1331 => x"06df3888",
  1332 => x"15811b70",
  1333 => x"8306555b",
  1334 => x"5572c938",
  1335 => x"7c830653",
  1336 => x"72802efd",
  1337 => x"b838ff1d",
  1338 => x"f819595d",
  1339 => x"88180878",
  1340 => x"2eea38fd",
  1341 => x"b539831a",
  1342 => x"53fc9639",
  1343 => x"83147082",
  1344 => x"2c81712b",
  1345 => x"80d7f808",
  1346 => x"077080d7",
  1347 => x"f40b8405",
  1348 => x"0c761010",
  1349 => x"1080d7f4",
  1350 => x"05881108",
  1351 => x"595b5e51",
  1352 => x"53fee139",
  1353 => x"80d7b808",
  1354 => x"1758b008",
  1355 => x"762e818d",
  1356 => x"3880d7e8",
  1357 => x"08ff2e83",
  1358 => x"ec387376",
  1359 => x"311880d7",
  1360 => x"b80c7387",
  1361 => x"06705753",
  1362 => x"72802e88",
  1363 => x"38887331",
  1364 => x"70155556",
  1365 => x"76149fff",
  1366 => x"06a08071",
  1367 => x"31177054",
  1368 => x"7f535753",
  1369 => x"84ee3fb0",
  1370 => x"0853b008",
  1371 => x"ff2e81a0",
  1372 => x"3880d7b8",
  1373 => x"08167080",
  1374 => x"d7b80c74",
  1375 => x"7580d7f4",
  1376 => x"0b88050c",
  1377 => x"74763118",
  1378 => x"70810751",
  1379 => x"5556587b",
  1380 => x"80d7f42e",
  1381 => x"839c3879",
  1382 => x"8f2682cb",
  1383 => x"38810b84",
  1384 => x"150c8415",
  1385 => x"08fc0670",
  1386 => x"7a317a72",
  1387 => x"268f7225",
  1388 => x"07525553",
  1389 => x"72802efc",
  1390 => x"f93880db",
  1391 => x"39b0089f",
  1392 => x"ff065372",
  1393 => x"feeb3877",
  1394 => x"80d7b80c",
  1395 => x"80d7f40b",
  1396 => x"8805087b",
  1397 => x"18810784",
  1398 => x"120c5580",
  1399 => x"d7e40878",
  1400 => x"27863877",
  1401 => x"80d7e40c",
  1402 => x"80d7e008",
  1403 => x"7827fcac",
  1404 => x"387780d7",
  1405 => x"e00c8415",
  1406 => x"08fc0670",
  1407 => x"7a317a72",
  1408 => x"268f7225",
  1409 => x"07525553",
  1410 => x"72802efc",
  1411 => x"a5388839",
  1412 => x"80745456",
  1413 => x"fedb397d",
  1414 => x"5183b83f",
  1415 => x"800bb00c",
  1416 => x"8f3d0d04",
  1417 => x"73538074",
  1418 => x"24a93872",
  1419 => x"822c8171",
  1420 => x"2b80d7f8",
  1421 => x"08077080",
  1422 => x"d7f40b84",
  1423 => x"050c5d53",
  1424 => x"778c180c",
  1425 => x"7488180c",
  1426 => x"7688190c",
  1427 => x"768c160c",
  1428 => x"f9b73983",
  1429 => x"1470822c",
  1430 => x"81712b80",
  1431 => x"d7f80807",
  1432 => x"7080d7f4",
  1433 => x"0b84050c",
  1434 => x"5e5153d4",
  1435 => x"397b7b06",
  1436 => x"5372fca3",
  1437 => x"38841a7b",
  1438 => x"105c5af1",
  1439 => x"39ff1a81",
  1440 => x"11515af7",
  1441 => x"b9397817",
  1442 => x"79810784",
  1443 => x"190c8c18",
  1444 => x"08881908",
  1445 => x"718c120c",
  1446 => x"88120c59",
  1447 => x"7080d888",
  1448 => x"0c7080d8",
  1449 => x"840c80d7",
  1450 => x"fc0b8c12",
  1451 => x"0c8c1108",
  1452 => x"88120c74",
  1453 => x"81078412",
  1454 => x"0c741175",
  1455 => x"710c5153",
  1456 => x"f9bd3975",
  1457 => x"17841108",
  1458 => x"81078412",
  1459 => x"0c538c17",
  1460 => x"08881808",
  1461 => x"718c120c",
  1462 => x"88120c58",
  1463 => x"7d5181f3",
  1464 => x"3f881754",
  1465 => x"f5cf3972",
  1466 => x"84150cf4",
  1467 => x"1af80670",
  1468 => x"841e0881",
  1469 => x"0607841e",
  1470 => x"0c701d54",
  1471 => x"5b850b84",
  1472 => x"140c850b",
  1473 => x"88140c8f",
  1474 => x"7b27fdcf",
  1475 => x"38881c52",
  1476 => x"7d518489",
  1477 => x"3f80d7f4",
  1478 => x"0b880508",
  1479 => x"80d7b808",
  1480 => x"5955fdb7",
  1481 => x"397780d7",
  1482 => x"b80c7380",
  1483 => x"d7e80cfc",
  1484 => x"91397284",
  1485 => x"150cfda3",
  1486 => x"39fc3d0d",
  1487 => x"7670797b",
  1488 => x"55555555",
  1489 => x"8f72278c",
  1490 => x"38727507",
  1491 => x"83065170",
  1492 => x"802ea738",
  1493 => x"ff125271",
  1494 => x"ff2e9838",
  1495 => x"72708105",
  1496 => x"54337470",
  1497 => x"81055634",
  1498 => x"ff125271",
  1499 => x"ff2e0981",
  1500 => x"06ea3874",
  1501 => x"b00c863d",
  1502 => x"0d047451",
  1503 => x"72708405",
  1504 => x"54087170",
  1505 => x"8405530c",
  1506 => x"72708405",
  1507 => x"54087170",
  1508 => x"8405530c",
  1509 => x"72708405",
  1510 => x"54087170",
  1511 => x"8405530c",
  1512 => x"72708405",
  1513 => x"54087170",
  1514 => x"8405530c",
  1515 => x"f0125271",
  1516 => x"8f26c938",
  1517 => x"83722795",
  1518 => x"38727084",
  1519 => x"05540871",
  1520 => x"70840553",
  1521 => x"0cfc1252",
  1522 => x"718326ed",
  1523 => x"387054ff",
  1524 => x"83390404",
  1525 => x"fd3d0d80",
  1526 => x"0b80e8c4",
  1527 => x"0c765189",
  1528 => x"d03fb008",
  1529 => x"53b008ff",
  1530 => x"2e883872",
  1531 => x"b00c853d",
  1532 => x"0d0480e8",
  1533 => x"c4085473",
  1534 => x"802ef038",
  1535 => x"7574710c",
  1536 => x"5272b00c",
  1537 => x"853d0d04",
  1538 => x"fd3d0d75",
  1539 => x"70718306",
  1540 => x"53555270",
  1541 => x"b8387170",
  1542 => x"087009f7",
  1543 => x"fbfdff12",
  1544 => x"0670f884",
  1545 => x"82818006",
  1546 => x"51515253",
  1547 => x"709d3884",
  1548 => x"13700870",
  1549 => x"09f7fbfd",
  1550 => x"ff120670",
  1551 => x"f8848281",
  1552 => x"80065151",
  1553 => x"52537080",
  1554 => x"2ee53872",
  1555 => x"52713351",
  1556 => x"70802e8a",
  1557 => x"38811270",
  1558 => x"33525270",
  1559 => x"f8387174",
  1560 => x"31b00c85",
  1561 => x"3d0d04fb",
  1562 => x"3d0d7770",
  1563 => x"5256fee2",
  1564 => x"3f80d7f4",
  1565 => x"0b880508",
  1566 => x"841108fc",
  1567 => x"06707b31",
  1568 => x"9fef05e0",
  1569 => x"8006e080",
  1570 => x"05565653",
  1571 => x"a0807424",
  1572 => x"94388052",
  1573 => x"7551febc",
  1574 => x"3f80d7fc",
  1575 => x"08155372",
  1576 => x"b0082e8f",
  1577 => x"387551fe",
  1578 => x"aa3f8053",
  1579 => x"72b00c87",
  1580 => x"3d0d0473",
  1581 => x"30527551",
  1582 => x"fe9a3fb0",
  1583 => x"08ff2ea8",
  1584 => x"3880d7f4",
  1585 => x"0b880508",
  1586 => x"75753181",
  1587 => x"0784120c",
  1588 => x"5380d7b8",
  1589 => x"08743180",
  1590 => x"d7b80c75",
  1591 => x"51fdf43f",
  1592 => x"810bb00c",
  1593 => x"873d0d04",
  1594 => x"80527551",
  1595 => x"fde63f80",
  1596 => x"d7f40b88",
  1597 => x"0508b008",
  1598 => x"71315653",
  1599 => x"8f7525ff",
  1600 => x"a438b008",
  1601 => x"80d7e808",
  1602 => x"3180d7b8",
  1603 => x"0c748107",
  1604 => x"84140c75",
  1605 => x"51fdbc3f",
  1606 => x"8053ff90",
  1607 => x"39f63d0d",
  1608 => x"7c7e545b",
  1609 => x"72802e82",
  1610 => x"83387a51",
  1611 => x"fda43ff8",
  1612 => x"13841108",
  1613 => x"70fe0670",
  1614 => x"13841108",
  1615 => x"fc065d58",
  1616 => x"59545880",
  1617 => x"d7fc0875",
  1618 => x"2e82de38",
  1619 => x"7884160c",
  1620 => x"80738106",
  1621 => x"545a727a",
  1622 => x"2e81d538",
  1623 => x"78158411",
  1624 => x"08810651",
  1625 => x"5372a038",
  1626 => x"78175779",
  1627 => x"81e63888",
  1628 => x"15085372",
  1629 => x"80d7fc2e",
  1630 => x"82f9388c",
  1631 => x"1508708c",
  1632 => x"150c7388",
  1633 => x"120c5676",
  1634 => x"81078419",
  1635 => x"0c761877",
  1636 => x"710c5379",
  1637 => x"81913883",
  1638 => x"ff772781",
  1639 => x"c8387689",
  1640 => x"2a77832a",
  1641 => x"56537280",
  1642 => x"2ebf3876",
  1643 => x"862ab805",
  1644 => x"55847327",
  1645 => x"b43880db",
  1646 => x"13559473",
  1647 => x"27ab3876",
  1648 => x"8c2a80ee",
  1649 => x"055580d4",
  1650 => x"73279e38",
  1651 => x"768f2a80",
  1652 => x"f7055582",
  1653 => x"d4732791",
  1654 => x"3876922a",
  1655 => x"80fc0555",
  1656 => x"8ad47327",
  1657 => x"843880fe",
  1658 => x"55741010",
  1659 => x"1080d7f4",
  1660 => x"05881108",
  1661 => x"55567376",
  1662 => x"2e82b338",
  1663 => x"841408fc",
  1664 => x"06537673",
  1665 => x"278d3888",
  1666 => x"14085473",
  1667 => x"762e0981",
  1668 => x"06ea388c",
  1669 => x"1408708c",
  1670 => x"1a0c7488",
  1671 => x"1a0c7888",
  1672 => x"120c5677",
  1673 => x"8c150c7a",
  1674 => x"51fba83f",
  1675 => x"8c3d0d04",
  1676 => x"77087871",
  1677 => x"31597705",
  1678 => x"88190854",
  1679 => x"577280d7",
  1680 => x"fc2e80e0",
  1681 => x"388c1808",
  1682 => x"708c150c",
  1683 => x"7388120c",
  1684 => x"56fe8939",
  1685 => x"8815088c",
  1686 => x"1608708c",
  1687 => x"130c5788",
  1688 => x"170cfea3",
  1689 => x"3976832a",
  1690 => x"70545580",
  1691 => x"75248198",
  1692 => x"3872822c",
  1693 => x"81712b80",
  1694 => x"d7f80807",
  1695 => x"80d7f40b",
  1696 => x"84050c53",
  1697 => x"74101010",
  1698 => x"80d7f405",
  1699 => x"88110855",
  1700 => x"56758c19",
  1701 => x"0c738819",
  1702 => x"0c778817",
  1703 => x"0c778c15",
  1704 => x"0cff8439",
  1705 => x"815afdb4",
  1706 => x"39781773",
  1707 => x"81065457",
  1708 => x"72983877",
  1709 => x"08787131",
  1710 => x"5977058c",
  1711 => x"1908881a",
  1712 => x"08718c12",
  1713 => x"0c88120c",
  1714 => x"57577681",
  1715 => x"0784190c",
  1716 => x"7780d7f4",
  1717 => x"0b88050c",
  1718 => x"80d7f008",
  1719 => x"7726fec7",
  1720 => x"3880d7ec",
  1721 => x"08527a51",
  1722 => x"fafd3f7a",
  1723 => x"51f9e43f",
  1724 => x"feba3981",
  1725 => x"788c150c",
  1726 => x"7888150c",
  1727 => x"738c1a0c",
  1728 => x"73881a0c",
  1729 => x"5afd8039",
  1730 => x"83157082",
  1731 => x"2c81712b",
  1732 => x"80d7f808",
  1733 => x"0780d7f4",
  1734 => x"0b84050c",
  1735 => x"51537410",
  1736 => x"101080d7",
  1737 => x"f4058811",
  1738 => x"085556fe",
  1739 => x"e4397453",
  1740 => x"807524a7",
  1741 => x"3872822c",
  1742 => x"81712b80",
  1743 => x"d7f80807",
  1744 => x"80d7f40b",
  1745 => x"84050c53",
  1746 => x"758c190c",
  1747 => x"7388190c",
  1748 => x"7788170c",
  1749 => x"778c150c",
  1750 => x"fdcd3983",
  1751 => x"1570822c",
  1752 => x"81712b80",
  1753 => x"d7f80807",
  1754 => x"80d7f40b",
  1755 => x"84050c51",
  1756 => x"53d639fc",
  1757 => x"3d0d7678",
  1758 => x"70085555",
  1759 => x"55728c38",
  1760 => x"73527451",
  1761 => x"fb973f86",
  1762 => x"3d0d0472",
  1763 => x"527451e3",
  1764 => x"3f735274",
  1765 => x"51fb863f",
  1766 => x"863d0d04",
  1767 => x"fb3d0d77",
  1768 => x"557480df",
  1769 => x"fc082e80",
  1770 => x"dd3880cc",
  1771 => x"15085380",
  1772 => x"5672762e",
  1773 => x"09810680",
  1774 => x"de3882c8",
  1775 => x"15085372",
  1776 => x"802ea338",
  1777 => x"82cc1556",
  1778 => x"72762e9a",
  1779 => x"38725475",
  1780 => x"742e9338",
  1781 => x"73740855",
  1782 => x"527451fa",
  1783 => x"c03f7574",
  1784 => x"2e098106",
  1785 => x"ef3880d4",
  1786 => x"15085372",
  1787 => x"80c238b8",
  1788 => x"1508802e",
  1789 => x"91387451",
  1790 => x"bc150853",
  1791 => x"722d84dc",
  1792 => x"15085372",
  1793 => x"b538873d",
  1794 => x"0d048116",
  1795 => x"56758e24",
  1796 => x"b43880cc",
  1797 => x"15085375",
  1798 => x"10101370",
  1799 => x"08555373",
  1800 => x"802ee738",
  1801 => x"73740855",
  1802 => x"527451f9",
  1803 => x"f03ff039",
  1804 => x"72527451",
  1805 => x"f9e73fff",
  1806 => x"b6397252",
  1807 => x"7451feb3",
  1808 => x"3f873d0d",
  1809 => x"0480cc15",
  1810 => x"08527451",
  1811 => x"f9cf3ffe",
  1812 => x"e939fb3d",
  1813 => x"0d775675",
  1814 => x"802e80c8",
  1815 => x"3882c816",
  1816 => x"08557480",
  1817 => x"2ea93884",
  1818 => x"1508ff05",
  1819 => x"54807424",
  1820 => x"98387310",
  1821 => x"10158805",
  1822 => x"537208fc",
  1823 => x"14545271",
  1824 => x"2dff1454",
  1825 => x"738025f1",
  1826 => x"38740855",
  1827 => x"74d938bc",
  1828 => x"16088538",
  1829 => x"873d0d04",
  1830 => x"7551bc16",
  1831 => x"0852712d",
  1832 => x"873d0d04",
  1833 => x"80dffc08",
  1834 => x"82c81108",
  1835 => x"5656ffb2",
  1836 => x"39fe3d0d",
  1837 => x"80e7fc08",
  1838 => x"51708a38",
  1839 => x"80e8c870",
  1840 => x"80e7fc0c",
  1841 => x"51707512",
  1842 => x"5252ff53",
  1843 => x"7087fb80",
  1844 => x"80268838",
  1845 => x"7080e7fc",
  1846 => x"0c715372",
  1847 => x"b00c843d",
  1848 => x"0d04fd3d",
  1849 => x"0d800b80",
  1850 => x"c9a80854",
  1851 => x"5472812e",
  1852 => x"9b387380",
  1853 => x"e8800ccf",
  1854 => x"ec3fce84",
  1855 => x"3f80e6fc",
  1856 => x"528151d2",
  1857 => x"8e3fb008",
  1858 => x"51879b3f",
  1859 => x"7280e880",
  1860 => x"0ccfd23f",
  1861 => x"cdea3f80",
  1862 => x"e6fc5281",
  1863 => x"51d1f43f",
  1864 => x"b0085187",
  1865 => x"813f00ff",
  1866 => x"3900ff39",
  1867 => x"f53d0d7e",
  1868 => x"6080e880",
  1869 => x"08705b58",
  1870 => x"5b5b7580",
  1871 => x"c238777a",
  1872 => x"25a13877",
  1873 => x"1b703370",
  1874 => x"81ff0658",
  1875 => x"5859758a",
  1876 => x"2e983876",
  1877 => x"81ff0651",
  1878 => x"ceea3f81",
  1879 => x"18587978",
  1880 => x"24e13879",
  1881 => x"b00c8d3d",
  1882 => x"0d048d51",
  1883 => x"ced63f78",
  1884 => x"337081ff",
  1885 => x"065257ce",
  1886 => x"cb3f8118",
  1887 => x"58e03979",
  1888 => x"557a547d",
  1889 => x"5385528d",
  1890 => x"3dfc0551",
  1891 => x"cdb33fb0",
  1892 => x"0856868b",
  1893 => x"3f7bb008",
  1894 => x"0c75b00c",
  1895 => x"8d3d0d04",
  1896 => x"f63d0d7d",
  1897 => x"7f80e880",
  1898 => x"08705b58",
  1899 => x"5a5a7580",
  1900 => x"c1387779",
  1901 => x"25b338cd",
  1902 => x"e63fb008",
  1903 => x"81ff0670",
  1904 => x"8d327030",
  1905 => x"709f2a51",
  1906 => x"51575776",
  1907 => x"8a2e80c3",
  1908 => x"3875802e",
  1909 => x"be38771a",
  1910 => x"56767634",
  1911 => x"7651cde4",
  1912 => x"3f811858",
  1913 => x"787824cf",
  1914 => x"38775675",
  1915 => x"b00c8c3d",
  1916 => x"0d047855",
  1917 => x"79547c53",
  1918 => x"84528c3d",
  1919 => x"fc0551cc",
  1920 => x"c03fb008",
  1921 => x"5685983f",
  1922 => x"7ab0080c",
  1923 => x"75b00c8c",
  1924 => x"3d0d0477",
  1925 => x"1a568a76",
  1926 => x"34811858",
  1927 => x"8d51cda4",
  1928 => x"3f8a51cd",
  1929 => x"9f3f7756",
  1930 => x"c239f93d",
  1931 => x"0d795780",
  1932 => x"e8800880",
  1933 => x"2eac3876",
  1934 => x"51f3cd3f",
  1935 => x"7b567a55",
  1936 => x"b0088105",
  1937 => x"54765382",
  1938 => x"52893dfc",
  1939 => x"0551cbf1",
  1940 => x"3fb00857",
  1941 => x"84c93f77",
  1942 => x"b0080c76",
  1943 => x"b00c893d",
  1944 => x"0d0484bb",
  1945 => x"3f850bb0",
  1946 => x"080cff0b",
  1947 => x"b00c893d",
  1948 => x"0d04fb3d",
  1949 => x"0d80e880",
  1950 => x"08705654",
  1951 => x"73883874",
  1952 => x"b00c873d",
  1953 => x"0d047753",
  1954 => x"8352873d",
  1955 => x"fc0551cb",
  1956 => x"b03fb008",
  1957 => x"5484883f",
  1958 => x"75b0080c",
  1959 => x"73b00c87",
  1960 => x"3d0d04ff",
  1961 => x"0bb00c04",
  1962 => x"fb3d0d77",
  1963 => x"5580e880",
  1964 => x"08802ea8",
  1965 => x"387451f2",
  1966 => x"cf3fb008",
  1967 => x"81055474",
  1968 => x"53875287",
  1969 => x"3dfc0551",
  1970 => x"caf73fb0",
  1971 => x"085583cf",
  1972 => x"3f75b008",
  1973 => x"0c74b00c",
  1974 => x"873d0d04",
  1975 => x"83c13f85",
  1976 => x"0bb0080c",
  1977 => x"ff0bb00c",
  1978 => x"873d0d04",
  1979 => x"fa3d0d80",
  1980 => x"e8800880",
  1981 => x"2ea2387a",
  1982 => x"55795478",
  1983 => x"53865288",
  1984 => x"3dfc0551",
  1985 => x"cabb3fb0",
  1986 => x"08568393",
  1987 => x"3f76b008",
  1988 => x"0c75b00c",
  1989 => x"883d0d04",
  1990 => x"83853f9d",
  1991 => x"0bb0080c",
  1992 => x"ff0bb00c",
  1993 => x"883d0d04",
  1994 => x"fb3d0d77",
  1995 => x"79565680",
  1996 => x"70545473",
  1997 => x"75259f38",
  1998 => x"74101010",
  1999 => x"f8055272",
  2000 => x"16703370",
  2001 => x"742b7607",
  2002 => x"8116f816",
  2003 => x"56565651",
  2004 => x"51747324",
  2005 => x"ea3873b0",
  2006 => x"0c873d0d",
  2007 => x"04fc3d0d",
  2008 => x"76785555",
  2009 => x"bc538052",
  2010 => x"735183de",
  2011 => x"3f845274",
  2012 => x"51ffb53f",
  2013 => x"b0087423",
  2014 => x"84528415",
  2015 => x"51ffa93f",
  2016 => x"b0088215",
  2017 => x"23845288",
  2018 => x"1551ff9c",
  2019 => x"3fb00884",
  2020 => x"150c8452",
  2021 => x"8c1551ff",
  2022 => x"8f3fb008",
  2023 => x"88152384",
  2024 => x"52901551",
  2025 => x"ff823fb0",
  2026 => x"088a1523",
  2027 => x"84529415",
  2028 => x"51fef53f",
  2029 => x"b0088c15",
  2030 => x"23845298",
  2031 => x"1551fee8",
  2032 => x"3fb0088e",
  2033 => x"15238852",
  2034 => x"9c1551fe",
  2035 => x"db3fb008",
  2036 => x"90150c86",
  2037 => x"3d0d04e9",
  2038 => x"3d0d6a80",
  2039 => x"e8800857",
  2040 => x"57759338",
  2041 => x"80c0800b",
  2042 => x"84180c75",
  2043 => x"ac180c75",
  2044 => x"b00c993d",
  2045 => x"0d04893d",
  2046 => x"70556a54",
  2047 => x"558a5299",
  2048 => x"3dffbc05",
  2049 => x"51c8ba3f",
  2050 => x"b0087753",
  2051 => x"755256fe",
  2052 => x"cc3f818b",
  2053 => x"3f77b008",
  2054 => x"0c75b00c",
  2055 => x"993d0d04",
  2056 => x"e93d0d69",
  2057 => x"5780e880",
  2058 => x"08802eb5",
  2059 => x"387651ef",
  2060 => x"d73f893d",
  2061 => x"7056b008",
  2062 => x"81055577",
  2063 => x"54568f52",
  2064 => x"993dffbc",
  2065 => x"0551c7f9",
  2066 => x"3fb0086b",
  2067 => x"53765257",
  2068 => x"fe8b3f80",
  2069 => x"ca3f77b0",
  2070 => x"080c76b0",
  2071 => x"0c993d0d",
  2072 => x"04bd3f85",
  2073 => x"0bb0080c",
  2074 => x"ff0bb00c",
  2075 => x"993d0d04",
  2076 => x"fc3d0d81",
  2077 => x"5480e880",
  2078 => x"08883873",
  2079 => x"b00c863d",
  2080 => x"0d047653",
  2081 => x"97b95286",
  2082 => x"3dfc0551",
  2083 => x"c7b33fb0",
  2084 => x"08548c3f",
  2085 => x"74b0080c",
  2086 => x"73b00c86",
  2087 => x"3d0d0480",
  2088 => x"dffc08b0",
  2089 => x"0c04f73d",
  2090 => x"0d7b80df",
  2091 => x"fc0882c8",
  2092 => x"11085a54",
  2093 => x"5a77802e",
  2094 => x"80da3881",
  2095 => x"88188419",
  2096 => x"08ff0581",
  2097 => x"712b5955",
  2098 => x"59807424",
  2099 => x"80ea3880",
  2100 => x"7424b538",
  2101 => x"73822b78",
  2102 => x"11880556",
  2103 => x"56818019",
  2104 => x"08770653",
  2105 => x"72802eb6",
  2106 => x"38781670",
  2107 => x"08535379",
  2108 => x"51740853",
  2109 => x"722dff14",
  2110 => x"fc17fc17",
  2111 => x"79812c5a",
  2112 => x"57575473",
  2113 => x"8025d638",
  2114 => x"77085877",
  2115 => x"ffad3880",
  2116 => x"dffc0853",
  2117 => x"bc1308a5",
  2118 => x"387951f8",
  2119 => x"893f7408",
  2120 => x"53722dff",
  2121 => x"14fc17fc",
  2122 => x"1779812c",
  2123 => x"5a575754",
  2124 => x"738025ff",
  2125 => x"a838d139",
  2126 => x"8057ff93",
  2127 => x"397251bc",
  2128 => x"13085372",
  2129 => x"2d7951f7",
  2130 => x"dd3ffc3d",
  2131 => x"0d767971",
  2132 => x"028c059f",
  2133 => x"05335755",
  2134 => x"53558372",
  2135 => x"278a3874",
  2136 => x"83065170",
  2137 => x"802ea238",
  2138 => x"ff125271",
  2139 => x"ff2e9338",
  2140 => x"73737081",
  2141 => x"055534ff",
  2142 => x"125271ff",
  2143 => x"2e098106",
  2144 => x"ef3874b0",
  2145 => x"0c863d0d",
  2146 => x"04747488",
  2147 => x"2b750770",
  2148 => x"71902b07",
  2149 => x"5154518f",
  2150 => x"7227a538",
  2151 => x"72717084",
  2152 => x"05530c72",
  2153 => x"71708405",
  2154 => x"530c7271",
  2155 => x"70840553",
  2156 => x"0c727170",
  2157 => x"8405530c",
  2158 => x"f0125271",
  2159 => x"8f26dd38",
  2160 => x"83722790",
  2161 => x"38727170",
  2162 => x"8405530c",
  2163 => x"fc125271",
  2164 => x"8326f238",
  2165 => x"7053ff90",
  2166 => x"39bc0802",
  2167 => x"bc0cfd3d",
  2168 => x"0d8053bc",
  2169 => x"088c0508",
  2170 => x"52bc0888",
  2171 => x"050851db",
  2172 => x"ff3fb008",
  2173 => x"70b00c54",
  2174 => x"853d0dbc",
  2175 => x"0c04bc08",
  2176 => x"02bc0cfd",
  2177 => x"3d0d8153",
  2178 => x"bc088c05",
  2179 => x"0852bc08",
  2180 => x"88050851",
  2181 => x"dbda3fb0",
  2182 => x"0870b00c",
  2183 => x"54853d0d",
  2184 => x"bc0c04ff",
  2185 => x"3d0d80e7",
  2186 => x"840bfc05",
  2187 => x"70085252",
  2188 => x"70ff2e91",
  2189 => x"38702dfc",
  2190 => x"12700852",
  2191 => x"5270ff2e",
  2192 => x"098106f1",
  2193 => x"38833d0d",
  2194 => x"0404c6e2",
  2195 => x"3f040000",
  2196 => x"00ffffff",
  2197 => x"ff00ffff",
  2198 => x"ffff00ff",
  2199 => x"ffffff00",
  2200 => x"00000040",
  2201 => x"75736167",
  2202 => x"653a2025",
  2203 => x"73202773",
  2204 => x"7472696e",
  2205 => x"67270a00",
  2206 => x"25322e32",
  2207 => x"78000000",
  2208 => x"00000007",
  2209 => x"0000000c",
  2210 => x"00000011",
  2211 => x"00000016",
  2212 => x"00000007",
  2213 => x"0000000c",
  2214 => x"00000011",
  2215 => x"00000016",
  2216 => x"00000007",
  2217 => x"0000000c",
  2218 => x"00000011",
  2219 => x"00000016",
  2220 => x"00000007",
  2221 => x"0000000c",
  2222 => x"00000011",
  2223 => x"00000016",
  2224 => x"00000005",
  2225 => x"00000009",
  2226 => x"0000000e",
  2227 => x"00000014",
  2228 => x"00000005",
  2229 => x"00000009",
  2230 => x"0000000e",
  2231 => x"00000014",
  2232 => x"00000005",
  2233 => x"00000009",
  2234 => x"0000000e",
  2235 => x"00000014",
  2236 => x"00000005",
  2237 => x"00000009",
  2238 => x"0000000e",
  2239 => x"00000014",
  2240 => x"00000004",
  2241 => x"0000000b",
  2242 => x"00000010",
  2243 => x"00000017",
  2244 => x"00000004",
  2245 => x"0000000b",
  2246 => x"00000010",
  2247 => x"00000017",
  2248 => x"00000004",
  2249 => x"0000000b",
  2250 => x"00000010",
  2251 => x"00000017",
  2252 => x"00000004",
  2253 => x"0000000b",
  2254 => x"00000010",
  2255 => x"00000017",
  2256 => x"00000006",
  2257 => x"0000000a",
  2258 => x"0000000f",
  2259 => x"00000015",
  2260 => x"00000006",
  2261 => x"0000000a",
  2262 => x"0000000f",
  2263 => x"00000015",
  2264 => x"00000006",
  2265 => x"0000000a",
  2266 => x"0000000f",
  2267 => x"00000015",
  2268 => x"00000006",
  2269 => x"0000000a",
  2270 => x"0000000f",
  2271 => x"00000015",
  2272 => x"d76aa478",
  2273 => x"e8c7b756",
  2274 => x"242070db",
  2275 => x"c1bdceee",
  2276 => x"f57c0faf",
  2277 => x"4787c62a",
  2278 => x"a8304613",
  2279 => x"fd469501",
  2280 => x"698098d8",
  2281 => x"8b44f7af",
  2282 => x"ffff5bb1",
  2283 => x"895cd7be",
  2284 => x"6b901122",
  2285 => x"fd987193",
  2286 => x"a679438e",
  2287 => x"49b40821",
  2288 => x"f61e2562",
  2289 => x"c040b340",
  2290 => x"265e5a51",
  2291 => x"e9b6c7aa",
  2292 => x"d62f105d",
  2293 => x"02441453",
  2294 => x"d8a1e681",
  2295 => x"e7d3fbc8",
  2296 => x"21e1cde6",
  2297 => x"c33707d6",
  2298 => x"f4d50d87",
  2299 => x"455a14ed",
  2300 => x"a9e3e905",
  2301 => x"fcefa3f8",
  2302 => x"676f02d9",
  2303 => x"8d2a4c8a",
  2304 => x"fffa3942",
  2305 => x"8771f681",
  2306 => x"6d9d6122",
  2307 => x"fde5380c",
  2308 => x"a4beea44",
  2309 => x"4bdecfa9",
  2310 => x"f6bb4b60",
  2311 => x"bebfbc70",
  2312 => x"289b7ec6",
  2313 => x"eaa127fa",
  2314 => x"d4ef3085",
  2315 => x"04881d05",
  2316 => x"d9d4d039",
  2317 => x"e6db99e5",
  2318 => x"1fa27cf8",
  2319 => x"c4ac5665",
  2320 => x"f4292244",
  2321 => x"432aff97",
  2322 => x"ab9423a7",
  2323 => x"fc93a039",
  2324 => x"655b59c3",
  2325 => x"8f0ccc92",
  2326 => x"ffeff47d",
  2327 => x"85845dd1",
  2328 => x"6fa87e4f",
  2329 => x"fe2ce6e0",
  2330 => x"a3014314",
  2331 => x"4e0811a1",
  2332 => x"f7537e82",
  2333 => x"bd3af235",
  2334 => x"2ad7d2bb",
  2335 => x"eb86d391",
  2336 => x"30313233",
  2337 => x"34353637",
  2338 => x"38394142",
  2339 => x"43444546",
  2340 => x"00000000",
  2341 => x"43000000",
  2342 => x"64756d6d",
  2343 => x"792e6578",
  2344 => x"65000000",
  2345 => x"00000000",
  2346 => x"00000000",
  2347 => x"00000000",
  2348 => x"0000338c",
  2349 => x"00000000",
  2350 => x"00000000",
  2351 => x"18181818",
  2352 => x"18001800",
  2353 => x"6c6c0000",
  2354 => x"00000000",
  2355 => x"6c6cfe6c",
  2356 => x"fe6c6c00",
  2357 => x"183e603c",
  2358 => x"067c1800",
  2359 => x"0066acd8",
  2360 => x"366acc00",
  2361 => x"386c6876",
  2362 => x"dcce7b00",
  2363 => x"18183000",
  2364 => x"00000000",
  2365 => x"0c183030",
  2366 => x"30180c00",
  2367 => x"30180c0c",
  2368 => x"0c183000",
  2369 => x"00663cff",
  2370 => x"3c660000",
  2371 => x"0018187e",
  2372 => x"18180000",
  2373 => x"00000000",
  2374 => x"00181830",
  2375 => x"0000007e",
  2376 => x"00000000",
  2377 => x"00000000",
  2378 => x"00181800",
  2379 => x"03060c18",
  2380 => x"3060c000",
  2381 => x"3c666e7e",
  2382 => x"76663c00",
  2383 => x"18387818",
  2384 => x"18181800",
  2385 => x"3c66060c",
  2386 => x"18307e00",
  2387 => x"3c66061c",
  2388 => x"06663c00",
  2389 => x"1c3c6ccc",
  2390 => x"fe0c0c00",
  2391 => x"7e607c06",
  2392 => x"06663c00",
  2393 => x"1c30607c",
  2394 => x"66663c00",
  2395 => x"7e06060c",
  2396 => x"18181800",
  2397 => x"3c66663c",
  2398 => x"66663c00",
  2399 => x"3c66663e",
  2400 => x"060c3800",
  2401 => x"00181800",
  2402 => x"00181800",
  2403 => x"00181800",
  2404 => x"00181830",
  2405 => x"00061860",
  2406 => x"18060000",
  2407 => x"00007e00",
  2408 => x"7e000000",
  2409 => x"00601806",
  2410 => x"18600000",
  2411 => x"3c66060c",
  2412 => x"18001800",
  2413 => x"7cc6ded6",
  2414 => x"dec07800",
  2415 => x"3c66667e",
  2416 => x"66666600",
  2417 => x"7c66667c",
  2418 => x"66667c00",
  2419 => x"1e306060",
  2420 => x"60301e00",
  2421 => x"786c6666",
  2422 => x"666c7800",
  2423 => x"7e606078",
  2424 => x"60607e00",
  2425 => x"7e606078",
  2426 => x"60606000",
  2427 => x"3c66606e",
  2428 => x"66663e00",
  2429 => x"6666667e",
  2430 => x"66666600",
  2431 => x"3c181818",
  2432 => x"18183c00",
  2433 => x"06060606",
  2434 => x"06663c00",
  2435 => x"c6ccd8f0",
  2436 => x"d8ccc600",
  2437 => x"60606060",
  2438 => x"60607e00",
  2439 => x"c6eefed6",
  2440 => x"c6c6c600",
  2441 => x"c6e6f6de",
  2442 => x"cec6c600",
  2443 => x"3c666666",
  2444 => x"66663c00",
  2445 => x"7c66667c",
  2446 => x"60606000",
  2447 => x"78cccccc",
  2448 => x"ccdc7e00",
  2449 => x"7c66667c",
  2450 => x"6c666600",
  2451 => x"3c66703c",
  2452 => x"0e663c00",
  2453 => x"7e181818",
  2454 => x"18181800",
  2455 => x"66666666",
  2456 => x"66663c00",
  2457 => x"66666666",
  2458 => x"3c3c1800",
  2459 => x"c6c6c6d6",
  2460 => x"feeec600",
  2461 => x"c3663c18",
  2462 => x"3c66c300",
  2463 => x"c3663c18",
  2464 => x"18181800",
  2465 => x"fe0c1830",
  2466 => x"60c0fe00",
  2467 => x"3c303030",
  2468 => x"30303c00",
  2469 => x"c0603018",
  2470 => x"0c060300",
  2471 => x"3c0c0c0c",
  2472 => x"0c0c3c00",
  2473 => x"10386cc6",
  2474 => x"00000000",
  2475 => x"00000000",
  2476 => x"000000fe",
  2477 => x"18180c00",
  2478 => x"00000000",
  2479 => x"00003c06",
  2480 => x"3e663e00",
  2481 => x"60607c66",
  2482 => x"66667c00",
  2483 => x"00003c60",
  2484 => x"60603c00",
  2485 => x"06063e66",
  2486 => x"66663e00",
  2487 => x"00003c66",
  2488 => x"7e603c00",
  2489 => x"1c307c30",
  2490 => x"30303000",
  2491 => x"00003e66",
  2492 => x"663e063c",
  2493 => x"60607c66",
  2494 => x"66666600",
  2495 => x"18001818",
  2496 => x"18180c00",
  2497 => x"0c000c0c",
  2498 => x"0c0c0c78",
  2499 => x"6060666c",
  2500 => x"786c6600",
  2501 => x"18181818",
  2502 => x"18180c00",
  2503 => x"0000ecfe",
  2504 => x"d6c6c600",
  2505 => x"00007c66",
  2506 => x"66666600",
  2507 => x"00003c66",
  2508 => x"66663c00",
  2509 => x"00007c66",
  2510 => x"667c6060",
  2511 => x"00003e66",
  2512 => x"663e0606",
  2513 => x"00007c66",
  2514 => x"60606000",
  2515 => x"00003c60",
  2516 => x"3c067c00",
  2517 => x"30307c30",
  2518 => x"30301c00",
  2519 => x"00006666",
  2520 => x"66663e00",
  2521 => x"00006666",
  2522 => x"663c1800",
  2523 => x"0000c6c6",
  2524 => x"d6fe6c00",
  2525 => x"0000c66c",
  2526 => x"386cc600",
  2527 => x"00006666",
  2528 => x"663c1830",
  2529 => x"00007e0c",
  2530 => x"18307e00",
  2531 => x"0e181870",
  2532 => x"18180e00",
  2533 => x"18181818",
  2534 => x"18181800",
  2535 => x"7018180e",
  2536 => x"18187000",
  2537 => x"729c0000",
  2538 => x"00000000",
  2539 => x"fefefefe",
  2540 => x"fefefe00",
  2541 => x"00000000",
  2542 => x"00000000",
  2543 => x"00000000",
  2544 => x"00000000",
  2545 => x"00000000",
  2546 => x"00000000",
  2547 => x"00000000",
  2548 => x"00000000",
  2549 => x"00000000",
  2550 => x"00000000",
  2551 => x"00000000",
  2552 => x"00000000",
  2553 => x"00000000",
  2554 => x"00000000",
  2555 => x"00000000",
  2556 => x"00000000",
  2557 => x"00000000",
  2558 => x"00000000",
  2559 => x"00000000",
  2560 => x"00000000",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"00000000",
  2564 => x"00000000",
  2565 => x"00000000",
  2566 => x"00000000",
  2567 => x"00000000",
  2568 => x"00000000",
  2569 => x"00000000",
  2570 => x"00000000",
  2571 => x"00000000",
  2572 => x"00000000",
  2573 => x"00000000",
  2574 => x"00000000",
  2575 => x"00000000",
  2576 => x"00000000",
  2577 => x"00000000",
  2578 => x"00000000",
  2579 => x"00000000",
  2580 => x"00000000",
  2581 => x"00000000",
  2582 => x"00000000",
  2583 => x"00000000",
  2584 => x"00000000",
  2585 => x"00000000",
  2586 => x"00000000",
  2587 => x"00000000",
  2588 => x"00000000",
  2589 => x"00000000",
  2590 => x"00000000",
  2591 => x"00000000",
  2592 => x"00000000",
  2593 => x"00000000",
  2594 => x"00000000",
  2595 => x"00000000",
  2596 => x"00000000",
  2597 => x"00000000",
  2598 => x"00000000",
  2599 => x"00000000",
  2600 => x"00000000",
  2601 => x"00000000",
  2602 => x"00000000",
  2603 => x"00000000",
  2604 => x"00000000",
  2605 => x"00000000",
  2606 => x"00000000",
  2607 => x"00000000",
  2608 => x"00000000",
  2609 => x"00000000",
  2610 => x"00000000",
  2611 => x"00000000",
  2612 => x"00000000",
  2613 => x"00000000",
  2614 => x"00000000",
  2615 => x"00000000",
  2616 => x"00000000",
  2617 => x"00000000",
  2618 => x"00000000",
  2619 => x"00000000",
  2620 => x"00000000",
  2621 => x"00000000",
  2622 => x"00000000",
  2623 => x"00000000",
  2624 => x"00000000",
  2625 => x"00000000",
  2626 => x"00000000",
  2627 => x"00000000",
  2628 => x"00000000",
  2629 => x"00000000",
  2630 => x"00000000",
  2631 => x"00000000",
  2632 => x"00000000",
  2633 => x"00000000",
  2634 => x"00000000",
  2635 => x"00000000",
  2636 => x"00000000",
  2637 => x"00000000",
  2638 => x"00000000",
  2639 => x"00000000",
  2640 => x"00000000",
  2641 => x"00000000",
  2642 => x"00000000",
  2643 => x"00000000",
  2644 => x"00000000",
  2645 => x"00000000",
  2646 => x"00000000",
  2647 => x"00000000",
  2648 => x"00000000",
  2649 => x"00000000",
  2650 => x"00000000",
  2651 => x"00000000",
  2652 => x"00000000",
  2653 => x"00000000",
  2654 => x"00000000",
  2655 => x"00000000",
  2656 => x"00000000",
  2657 => x"00000000",
  2658 => x"00000000",
  2659 => x"00000000",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000000",
  2683 => x"00000000",
  2684 => x"00000000",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000000",
  2712 => x"00000000",
  2713 => x"00000000",
  2714 => x"00000000",
  2715 => x"00000000",
  2716 => x"00000000",
  2717 => x"00000000",
  2718 => x"00000000",
  2719 => x"00000000",
  2720 => x"00000000",
  2721 => x"00000000",
  2722 => x"00000000",
  2723 => x"00000000",
  2724 => x"00000000",
  2725 => x"00000000",
  2726 => x"00000000",
  2727 => x"00000000",
  2728 => x"00000000",
  2729 => x"00000000",
  2730 => x"00000000",
  2731 => x"00000000",
  2732 => x"00000000",
  2733 => x"00000000",
  2734 => x"00000000",
  2735 => x"00000000",
  2736 => x"00000000",
  2737 => x"00000000",
  2738 => x"00000000",
  2739 => x"00000000",
  2740 => x"00000000",
  2741 => x"00000000",
  2742 => x"00000000",
  2743 => x"00000000",
  2744 => x"00000000",
  2745 => x"00000000",
  2746 => x"00000000",
  2747 => x"00000000",
  2748 => x"00000000",
  2749 => x"00000000",
  2750 => x"00000000",
  2751 => x"00000000",
  2752 => x"00000000",
  2753 => x"00000000",
  2754 => x"00000000",
  2755 => x"00000000",
  2756 => x"00000000",
  2757 => x"00000000",
  2758 => x"00000000",
  2759 => x"00000000",
  2760 => x"00000000",
  2761 => x"00000000",
  2762 => x"00000000",
  2763 => x"00000000",
  2764 => x"00000000",
  2765 => x"00000000",
  2766 => x"00000000",
  2767 => x"00000000",
  2768 => x"00000000",
  2769 => x"00000000",
  2770 => x"00000000",
  2771 => x"00000000",
  2772 => x"00000000",
  2773 => x"00000000",
  2774 => x"00000000",
  2775 => x"00000000",
  2776 => x"00000000",
  2777 => x"00000000",
  2778 => x"00000000",
  2779 => x"00000000",
  2780 => x"00000000",
  2781 => x"00000000",
  2782 => x"00000000",
  2783 => x"00000000",
  2784 => x"00000000",
  2785 => x"00000000",
  2786 => x"00000000",
  2787 => x"00000000",
  2788 => x"00000000",
  2789 => x"00000000",
  2790 => x"00000000",
  2791 => x"00000000",
  2792 => x"00000000",
  2793 => x"00000000",
  2794 => x"00000000",
  2795 => x"00000000",
  2796 => x"00000000",
  2797 => x"0000c100",
  2798 => x"00000000",
  2799 => x"00000000",
  2800 => x"00000000",
  2801 => x"00000000",
  2802 => x"00000000",
  2803 => x"00000000",
  2804 => x"00000000",
  2805 => x"00000000",
  2806 => x"00000000",
  2807 => x"00000000",
  2808 => x"00000000",
  2809 => x"00000000",
  2810 => x"ffffffff",
  2811 => x"00000000",
  2812 => x"00020000",
  2813 => x"00000000",
  2814 => x"00000000",
  2815 => x"00002bf4",
  2816 => x"00002bf4",
  2817 => x"00002bfc",
  2818 => x"00002bfc",
  2819 => x"00002c04",
  2820 => x"00002c04",
  2821 => x"00002c0c",
  2822 => x"00002c0c",
  2823 => x"00002c14",
  2824 => x"00002c14",
  2825 => x"00002c1c",
  2826 => x"00002c1c",
  2827 => x"00002c24",
  2828 => x"00002c24",
  2829 => x"00002c2c",
  2830 => x"00002c2c",
  2831 => x"00002c34",
  2832 => x"00002c34",
  2833 => x"00002c3c",
  2834 => x"00002c3c",
  2835 => x"00002c44",
  2836 => x"00002c44",
  2837 => x"00002c4c",
  2838 => x"00002c4c",
  2839 => x"00002c54",
  2840 => x"00002c54",
  2841 => x"00002c5c",
  2842 => x"00002c5c",
  2843 => x"00002c64",
  2844 => x"00002c64",
  2845 => x"00002c6c",
  2846 => x"00002c6c",
  2847 => x"00002c74",
  2848 => x"00002c74",
  2849 => x"00002c7c",
  2850 => x"00002c7c",
  2851 => x"00002c84",
  2852 => x"00002c84",
  2853 => x"00002c8c",
  2854 => x"00002c8c",
  2855 => x"00002c94",
  2856 => x"00002c94",
  2857 => x"00002c9c",
  2858 => x"00002c9c",
  2859 => x"00002ca4",
  2860 => x"00002ca4",
  2861 => x"00002cac",
  2862 => x"00002cac",
  2863 => x"00002cb4",
  2864 => x"00002cb4",
  2865 => x"00002cbc",
  2866 => x"00002cbc",
  2867 => x"00002cc4",
  2868 => x"00002cc4",
  2869 => x"00002ccc",
  2870 => x"00002ccc",
  2871 => x"00002cd4",
  2872 => x"00002cd4",
  2873 => x"00002cdc",
  2874 => x"00002cdc",
  2875 => x"00002ce4",
  2876 => x"00002ce4",
  2877 => x"00002cec",
  2878 => x"00002cec",
  2879 => x"00002cf4",
  2880 => x"00002cf4",
  2881 => x"00002cfc",
  2882 => x"00002cfc",
  2883 => x"00002d04",
  2884 => x"00002d04",
  2885 => x"00002d0c",
  2886 => x"00002d0c",
  2887 => x"00002d14",
  2888 => x"00002d14",
  2889 => x"00002d1c",
  2890 => x"00002d1c",
  2891 => x"00002d24",
  2892 => x"00002d24",
  2893 => x"00002d2c",
  2894 => x"00002d2c",
  2895 => x"00002d34",
  2896 => x"00002d34",
  2897 => x"00002d3c",
  2898 => x"00002d3c",
  2899 => x"00002d44",
  2900 => x"00002d44",
  2901 => x"00002d4c",
  2902 => x"00002d4c",
  2903 => x"00002d54",
  2904 => x"00002d54",
  2905 => x"00002d5c",
  2906 => x"00002d5c",
  2907 => x"00002d64",
  2908 => x"00002d64",
  2909 => x"00002d6c",
  2910 => x"00002d6c",
  2911 => x"00002d74",
  2912 => x"00002d74",
  2913 => x"00002d7c",
  2914 => x"00002d7c",
  2915 => x"00002d84",
  2916 => x"00002d84",
  2917 => x"00002d8c",
  2918 => x"00002d8c",
  2919 => x"00002d94",
  2920 => x"00002d94",
  2921 => x"00002d9c",
  2922 => x"00002d9c",
  2923 => x"00002da4",
  2924 => x"00002da4",
  2925 => x"00002dac",
  2926 => x"00002dac",
  2927 => x"00002db4",
  2928 => x"00002db4",
  2929 => x"00002dbc",
  2930 => x"00002dbc",
  2931 => x"00002dc4",
  2932 => x"00002dc4",
  2933 => x"00002dcc",
  2934 => x"00002dcc",
  2935 => x"00002dd4",
  2936 => x"00002dd4",
  2937 => x"00002ddc",
  2938 => x"00002ddc",
  2939 => x"00002de4",
  2940 => x"00002de4",
  2941 => x"00002dec",
  2942 => x"00002dec",
  2943 => x"00002df4",
  2944 => x"00002df4",
  2945 => x"00002dfc",
  2946 => x"00002dfc",
  2947 => x"00002e04",
  2948 => x"00002e04",
  2949 => x"00002e0c",
  2950 => x"00002e0c",
  2951 => x"00002e14",
  2952 => x"00002e14",
  2953 => x"00002e1c",
  2954 => x"00002e1c",
  2955 => x"00002e24",
  2956 => x"00002e24",
  2957 => x"00002e2c",
  2958 => x"00002e2c",
  2959 => x"00002e34",
  2960 => x"00002e34",
  2961 => x"00002e3c",
  2962 => x"00002e3c",
  2963 => x"00002e44",
  2964 => x"00002e44",
  2965 => x"00002e4c",
  2966 => x"00002e4c",
  2967 => x"00002e54",
  2968 => x"00002e54",
  2969 => x"00002e5c",
  2970 => x"00002e5c",
  2971 => x"00002e64",
  2972 => x"00002e64",
  2973 => x"00002e6c",
  2974 => x"00002e6c",
  2975 => x"00002e74",
  2976 => x"00002e74",
  2977 => x"00002e7c",
  2978 => x"00002e7c",
  2979 => x"00002e84",
  2980 => x"00002e84",
  2981 => x"00002e8c",
  2982 => x"00002e8c",
  2983 => x"00002e94",
  2984 => x"00002e94",
  2985 => x"00002e9c",
  2986 => x"00002e9c",
  2987 => x"00002ea4",
  2988 => x"00002ea4",
  2989 => x"00002eac",
  2990 => x"00002eac",
  2991 => x"00002eb4",
  2992 => x"00002eb4",
  2993 => x"00002ebc",
  2994 => x"00002ebc",
  2995 => x"00002ec4",
  2996 => x"00002ec4",
  2997 => x"00002ecc",
  2998 => x"00002ecc",
  2999 => x"00002ed4",
  3000 => x"00002ed4",
  3001 => x"00002edc",
  3002 => x"00002edc",
  3003 => x"00002ee4",
  3004 => x"00002ee4",
  3005 => x"00002eec",
  3006 => x"00002eec",
  3007 => x"00002ef4",
  3008 => x"00002ef4",
  3009 => x"00002efc",
  3010 => x"00002efc",
  3011 => x"00002f04",
  3012 => x"00002f04",
  3013 => x"00002f0c",
  3014 => x"00002f0c",
  3015 => x"00002f14",
  3016 => x"00002f14",
  3017 => x"00002f1c",
  3018 => x"00002f1c",
  3019 => x"00002f24",
  3020 => x"00002f24",
  3021 => x"00002f2c",
  3022 => x"00002f2c",
  3023 => x"00002f34",
  3024 => x"00002f34",
  3025 => x"00002f3c",
  3026 => x"00002f3c",
  3027 => x"00002f44",
  3028 => x"00002f44",
  3029 => x"00002f4c",
  3030 => x"00002f4c",
  3031 => x"00002f54",
  3032 => x"00002f54",
  3033 => x"00002f5c",
  3034 => x"00002f5c",
  3035 => x"00002f64",
  3036 => x"00002f64",
  3037 => x"00002f6c",
  3038 => x"00002f6c",
  3039 => x"00002f74",
  3040 => x"00002f74",
  3041 => x"00002f7c",
  3042 => x"00002f7c",
  3043 => x"00002f84",
  3044 => x"00002f84",
  3045 => x"00002f8c",
  3046 => x"00002f8c",
  3047 => x"00002f94",
  3048 => x"00002f94",
  3049 => x"00002f9c",
  3050 => x"00002f9c",
  3051 => x"00002fa4",
  3052 => x"00002fa4",
  3053 => x"00002fac",
  3054 => x"00002fac",
  3055 => x"00002fb4",
  3056 => x"00002fb4",
  3057 => x"00002fbc",
  3058 => x"00002fbc",
  3059 => x"00002fc4",
  3060 => x"00002fc4",
  3061 => x"00002fcc",
  3062 => x"00002fcc",
  3063 => x"00002fd4",
  3064 => x"00002fd4",
  3065 => x"00002fdc",
  3066 => x"00002fdc",
  3067 => x"00002fe4",
  3068 => x"00002fe4",
  3069 => x"00002fec",
  3070 => x"00002fec",
  3071 => x"00003000",
  3072 => x"00000000",
  3073 => x"00003268",
  3074 => x"000032c4",
  3075 => x"00003320",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000000",
  3084 => x"00000000",
  3085 => x"00002494",
  3086 => x"00000000",
  3087 => x"00000000",
  3088 => x"00000000",
  3089 => x"00000000",
  3090 => x"00000000",
  3091 => x"00000000",
  3092 => x"00000000",
  3093 => x"00000000",
  3094 => x"00000000",
  3095 => x"00000000",
  3096 => x"00000000",
  3097 => x"00000000",
  3098 => x"00000000",
  3099 => x"00000000",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00000000",
  3103 => x"00000000",
  3104 => x"00000000",
  3105 => x"00000000",
  3106 => x"00000000",
  3107 => x"00000000",
  3108 => x"00000000",
  3109 => x"00000000",
  3110 => x"00000000",
  3111 => x"00000000",
  3112 => x"00000000",
  3113 => x"00000000",
  3114 => x"00000001",
  3115 => x"330eabcd",
  3116 => x"1234e66d",
  3117 => x"deec0005",
  3118 => x"000b0000",
  3119 => x"00000000",
  3120 => x"00000000",
  3121 => x"00000000",
  3122 => x"00000000",
  3123 => x"00000000",
  3124 => x"00000000",
  3125 => x"00000000",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000000",
  3151 => x"00000000",
  3152 => x"00000000",
  3153 => x"00000000",
  3154 => x"00000000",
  3155 => x"00000000",
  3156 => x"00000000",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"00000000",
  3161 => x"00000000",
  3162 => x"00000000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"00000000",
  3166 => x"00000000",
  3167 => x"00000000",
  3168 => x"00000000",
  3169 => x"00000000",
  3170 => x"00000000",
  3171 => x"00000000",
  3172 => x"00000000",
  3173 => x"00000000",
  3174 => x"00000000",
  3175 => x"00000000",
  3176 => x"00000000",
  3177 => x"00000000",
  3178 => x"00000000",
  3179 => x"00000000",
  3180 => x"00000000",
  3181 => x"00000000",
  3182 => x"00000000",
  3183 => x"00000000",
  3184 => x"00000000",
  3185 => x"00000000",
  3186 => x"00000000",
  3187 => x"00000000",
  3188 => x"00000000",
  3189 => x"00000000",
  3190 => x"00000000",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00000000",
  3195 => x"00000000",
  3196 => x"00000000",
  3197 => x"00000000",
  3198 => x"00000000",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"00000000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000000",
  3246 => x"00000000",
  3247 => x"00000000",
  3248 => x"00000000",
  3249 => x"00000000",
  3250 => x"00000000",
  3251 => x"00000000",
  3252 => x"00000000",
  3253 => x"00000000",
  3254 => x"00000000",
  3255 => x"00000000",
  3256 => x"00000000",
  3257 => x"00000000",
  3258 => x"00000000",
  3259 => x"00000000",
  3260 => x"00000000",
  3261 => x"00000000",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00000000",
  3265 => x"00000000",
  3266 => x"00000000",
  3267 => x"00000000",
  3268 => x"00000000",
  3269 => x"00000000",
  3270 => x"00000000",
  3271 => x"00000000",
  3272 => x"00000000",
  3273 => x"00000000",
  3274 => x"00000000",
  3275 => x"00000000",
  3276 => x"00000000",
  3277 => x"00000000",
  3278 => x"00000000",
  3279 => x"00000000",
  3280 => x"00000000",
  3281 => x"00000000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"00000000",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00000000",
  3288 => x"00000000",
  3289 => x"00000000",
  3290 => x"00000000",
  3291 => x"00000000",
  3292 => x"00000000",
  3293 => x"00000000",
  3294 => x"00000000",
  3295 => x"00002498",
  3296 => x"ffffffff",
  3297 => x"00000000",
  3298 => x"ffffffff",
  3299 => x"00000000",
  3300 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

