-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a0808491",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"8bb87383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02ec050d",
    30 => x"76548755",
    31 => x"739c2a74",
    32 => x"842bb712",
    33 => x"55555271",
    34 => x"89248438",
    35 => x"b0125372",
    36 => x"51a08087",
    37 => x"ba2dff15",
    38 => x"55748025",
    39 => x"df380294",
    40 => x"050d0402",
    41 => x"e8050d87",
    42 => x"f0808008",
    43 => x"9e800a08",
    44 => x"55568755",
    45 => x"739c2a74",
    46 => x"842bb712",
    47 => x"55555271",
    48 => x"89248438",
    49 => x"b0125372",
    50 => x"51a08087",
    51 => x"ba2dff15",
    52 => x"55748025",
    53 => x"df387554",
    54 => x"8755739c",
    55 => x"2a74842b",
    56 => x"b7125555",
    57 => x"52718924",
    58 => x"8438b012",
    59 => x"537251a0",
    60 => x"8087ba2d",
    61 => x"ff155574",
    62 => x"8025df38",
    63 => x"87f08084",
    64 => x"0887c080",
    65 => x"84085556",
    66 => x"8755739c",
    67 => x"2a74842b",
    68 => x"b7125555",
    69 => x"52718924",
    70 => x"8438b012",
    71 => x"537251a0",
    72 => x"8087ba2d",
    73 => x"ff155574",
    74 => x"8025df38",
    75 => x"75548755",
    76 => x"739c2a74",
    77 => x"842bb712",
    78 => x"55555271",
    79 => x"89248438",
    80 => x"b0125372",
    81 => x"51a08087",
    82 => x"ba2dff15",
    83 => x"55748025",
    84 => x"df388a51",
    85 => x"a08087ba",
    86 => x"2d87f080",
    87 => x"880887c0",
    88 => x"80880855",
    89 => x"56875573",
    90 => x"9c2a7484",
    91 => x"2bb71255",
    92 => x"55527189",
    93 => x"248438b0",
    94 => x"12537251",
    95 => x"a08087ba",
    96 => x"2dff1555",
    97 => x"748025df",
    98 => x"38755487",
    99 => x"55739c2a",
   100 => x"74842bb7",
   101 => x"12555552",
   102 => x"71892484",
   103 => x"38b01253",
   104 => x"7251a080",
   105 => x"87ba2dff",
   106 => x"15557480",
   107 => x"25df3887",
   108 => x"f0808c08",
   109 => x"87c0808c",
   110 => x"08555687",
   111 => x"55739c2a",
   112 => x"74842bb7",
   113 => x"12555552",
   114 => x"71892484",
   115 => x"38b01253",
   116 => x"7251a080",
   117 => x"87ba2dff",
   118 => x"15557480",
   119 => x"25df3875",
   120 => x"54875573",
   121 => x"9c2a7484",
   122 => x"2bb71255",
   123 => x"55527189",
   124 => x"248438b0",
   125 => x"12537251",
   126 => x"a08087ba",
   127 => x"2dff1555",
   128 => x"748025df",
   129 => x"388a51a0",
   130 => x"8087ba2d",
   131 => x"0298050d",
   132 => x"0402f805",
   133 => x"0d830b85",
   134 => x"ffc48134",
   135 => x"fc0b85ff",
   136 => x"c08134a0",
   137 => x"8084f62d",
   138 => x"80c851a0",
   139 => x"8087ba2d",
   140 => x"80e551a0",
   141 => x"8087ba2d",
   142 => x"80ec51a0",
   143 => x"8087ba2d",
   144 => x"80ec51a0",
   145 => x"8087ba2d",
   146 => x"80ef51a0",
   147 => x"8087ba2d",
   148 => x"8a51a080",
   149 => x"87ba2da0",
   150 => x"808bc851",
   151 => x"a08089a1",
   152 => x"2d87f080",
   153 => x"8022529e",
   154 => x"800a229e",
   155 => x"800a2251",
   156 => x"52a08084",
   157 => x"e70402f4",
   158 => x"050dfea0",
   159 => x"800b86ff",
   160 => x"e2802380",
   161 => x"0b86ffe2",
   162 => x"8223800b",
   163 => x"86ffe284",
   164 => x"23800b86",
   165 => x"ffe28823",
   166 => x"800b86ff",
   167 => x"e28a2390",
   168 => x"705353a0",
   169 => x"bf518072",
   170 => x"70840554",
   171 => x"0cff1151",
   172 => x"708025f2",
   173 => x"38bc0b86",
   174 => x"ffe19223",
   175 => x"81d40b86",
   176 => x"ffe19423",
   177 => x"80d9810b",
   178 => x"86ffe18e",
   179 => x"23e9c10b",
   180 => x"86ffe190",
   181 => x"2386ff0b",
   182 => x"86ffe380",
   183 => x"239fff0b",
   184 => x"86ffe382",
   185 => x"2381e00b",
   186 => x"84889023",
   187 => x"900b902c",
   188 => x"51708488",
   189 => x"922381e2",
   190 => x"0b848894",
   191 => x"23728488",
   192 => x"9623ff0b",
   193 => x"84889823",
   194 => x"fe0b8488",
   195 => x"9a238488",
   196 => x"900b902c",
   197 => x"527186ff",
   198 => x"e1802384",
   199 => x"88905170",
   200 => x"86ffe182",
   201 => x"23800b86",
   202 => x"ffe18823",
   203 => x"fe87900b",
   204 => x"86ffe196",
   205 => x"23800b84",
   206 => x"88a00c80",
   207 => x"0b8488a4",
   208 => x"0c028c05",
   209 => x"0d0402f8",
   210 => x"050d8488",
   211 => x"a4081010",
   212 => x"8488a408",
   213 => x"05709029",
   214 => x"8488a008",
   215 => x"0584c011",
   216 => x"51525280",
   217 => x"52717134",
   218 => x"71811234",
   219 => x"71821234",
   220 => x"71831234",
   221 => x"80d01181",
   222 => x"13535181",
   223 => x"ff7225e5",
   224 => x"38028805",
   225 => x"0d0402f4",
   226 => x"050d9053",
   227 => x"a0bf5272",
   228 => x"84147108",
   229 => x"8105720c",
   230 => x"ff145454",
   231 => x"51807224",
   232 => x"e9387284",
   233 => x"14710881",
   234 => x"05720cff",
   235 => x"14545451",
   236 => x"718025db",
   237 => x"38a08087",
   238 => x"8a0402e8",
   239 => x"050d7756",
   240 => x"9f762581",
   241 => x"8d388488",
   242 => x"a4087010",
   243 => x"10117081",
   244 => x"80298488",
   245 => x"a0080584",
   246 => x"c0117910",
   247 => x"1010a080",
   248 => x"89d80570",
   249 => x"70840552",
   250 => x"08710852",
   251 => x"54555154",
   252 => x"55557072",
   253 => x"3470882c",
   254 => x"5372ffb0",
   255 => x"13347090",
   256 => x"2c5372fe",
   257 => x"e0133470",
   258 => x"982c5170",
   259 => x"fe901334",
   260 => x"73fdc013",
   261 => x"3473882c",
   262 => x"5372fcf0",
   263 => x"13347390",
   264 => x"2c5170fc",
   265 => x"a0133473",
   266 => x"982c5473",
   267 => x"fbd01334",
   268 => x"758a2eab",
   269 => x"388488a0",
   270 => x"08810584",
   271 => x"88a00c84",
   272 => x"88a00880",
   273 => x"d02e9838",
   274 => x"74992eac",
   275 => x"38029805",
   276 => x"0d048488",
   277 => x"a4085575",
   278 => x"8a2e0981",
   279 => x"06d73881",
   280 => x"158488a4",
   281 => x"0c800b84",
   282 => x"88a00c84",
   283 => x"88a40855",
   284 => x"74992e09",
   285 => x"8106d638",
   286 => x"900b9480",
   287 => x"1154529f",
   288 => x"9f517270",
   289 => x"84055408",
   290 => x"72708405",
   291 => x"540cff11",
   292 => x"51708025",
   293 => x"ed38980b",
   294 => x"8488a40c",
   295 => x"0298050d",
   296 => x"0402dc05",
   297 => x"0d7a5877",
   298 => x"70840559",
   299 => x"08578059",
   300 => x"76982a77",
   301 => x"882b5856",
   302 => x"75802e81",
   303 => x"9b389f76",
   304 => x"25819a38",
   305 => x"8488a408",
   306 => x"70101011",
   307 => x"70818029",
   308 => x"8488a008",
   309 => x"0584c011",
   310 => x"79101010",
   311 => x"a08089d8",
   312 => x"05707084",
   313 => x"05520871",
   314 => x"08525455",
   315 => x"51545555",
   316 => x"70723470",
   317 => x"882c5372",
   318 => x"ffb01334",
   319 => x"70902c53",
   320 => x"72fee013",
   321 => x"3470982c",
   322 => x"5170fe90",
   323 => x"133473fd",
   324 => x"c0133473",
   325 => x"882c5372",
   326 => x"fcf01334",
   327 => x"73902c51",
   328 => x"70fca013",
   329 => x"3473982c",
   330 => x"5473fbd0",
   331 => x"1334758a",
   332 => x"2eb83884",
   333 => x"88a00881",
   334 => x"058488a0",
   335 => x"0c8488a0",
   336 => x"0880d02e",
   337 => x"a5387499",
   338 => x"2eb93881",
   339 => x"19598379",
   340 => x"25fedd38",
   341 => x"75fed038",
   342 => x"02a4050d",
   343 => x"048488a4",
   344 => x"0855758a",
   345 => x"2e098106",
   346 => x"ca388115",
   347 => x"8488a40c",
   348 => x"800b8488",
   349 => x"a00c8488",
   350 => x"a4085574",
   351 => x"992e0981",
   352 => x"06c93890",
   353 => x"0b948011",
   354 => x"54529f9f",
   355 => x"51727084",
   356 => x"05540872",
   357 => x"70840554",
   358 => x"0cff1151",
   359 => x"708025ed",
   360 => x"38980b84",
   361 => x"88a40c81",
   362 => x"19598379",
   363 => x"25fe8138",
   364 => x"a0808ad4",
   365 => x"04000000",
   366 => x"00ffffff",
   367 => x"ff00ffff",
   368 => x"ffff00ff",
   369 => x"ffffff00",
   370 => x"48656c6c",
   371 => x"6f2c2077",
   372 => x"6f726c64",
   373 => x"210a0000",
   374 => x"00000000",
   375 => x"00000000",
   376 => x"18181818",
   377 => x"18001800",
   378 => x"6c6c0000",
   379 => x"00000000",
   380 => x"6c6cfe6c",
   381 => x"fe6c6c00",
   382 => x"183e603c",
   383 => x"067c1800",
   384 => x"0066acd8",
   385 => x"366acc00",
   386 => x"386c6876",
   387 => x"dcce7b00",
   388 => x"18183000",
   389 => x"00000000",
   390 => x"0c183030",
   391 => x"30180c00",
   392 => x"30180c0c",
   393 => x"0c183000",
   394 => x"00663cff",
   395 => x"3c660000",
   396 => x"0018187e",
   397 => x"18180000",
   398 => x"00000000",
   399 => x"00181830",
   400 => x"0000007e",
   401 => x"00000000",
   402 => x"00000000",
   403 => x"00181800",
   404 => x"03060c18",
   405 => x"3060c000",
   406 => x"3c666e7e",
   407 => x"76663c00",
   408 => x"18387818",
   409 => x"18181800",
   410 => x"3c66060c",
   411 => x"18307e00",
   412 => x"3c66061c",
   413 => x"06663c00",
   414 => x"1c3c6ccc",
   415 => x"fe0c0c00",
   416 => x"7e607c06",
   417 => x"06663c00",
   418 => x"1c30607c",
   419 => x"66663c00",
   420 => x"7e06060c",
   421 => x"18181800",
   422 => x"3c66663c",
   423 => x"66663c00",
   424 => x"3c66663e",
   425 => x"060c3800",
   426 => x"00181800",
   427 => x"00181800",
   428 => x"00181800",
   429 => x"00181830",
   430 => x"00061860",
   431 => x"18060000",
   432 => x"00007e00",
   433 => x"7e000000",
   434 => x"00601806",
   435 => x"18600000",
   436 => x"3c66060c",
   437 => x"18001800",
   438 => x"7cc6ded6",
   439 => x"dec07800",
   440 => x"3c66667e",
   441 => x"66666600",
   442 => x"7c66667c",
   443 => x"66667c00",
   444 => x"1e306060",
   445 => x"60301e00",
   446 => x"786c6666",
   447 => x"666c7800",
   448 => x"7e606078",
   449 => x"60607e00",
   450 => x"7e606078",
   451 => x"60606000",
   452 => x"3c66606e",
   453 => x"66663e00",
   454 => x"6666667e",
   455 => x"66666600",
   456 => x"3c181818",
   457 => x"18183c00",
   458 => x"06060606",
   459 => x"06663c00",
   460 => x"c6ccd8f0",
   461 => x"d8ccc600",
   462 => x"60606060",
   463 => x"60607e00",
   464 => x"c6eefed6",
   465 => x"c6c6c600",
   466 => x"c6e6f6de",
   467 => x"cec6c600",
   468 => x"3c666666",
   469 => x"66663c00",
   470 => x"7c66667c",
   471 => x"60606000",
   472 => x"78cccccc",
   473 => x"ccdc7e00",
   474 => x"7c66667c",
   475 => x"6c666600",
   476 => x"3c66703c",
   477 => x"0e663c00",
   478 => x"7e181818",
   479 => x"18181800",
   480 => x"66666666",
   481 => x"66663c00",
   482 => x"66666666",
   483 => x"3c3c1800",
   484 => x"c6c6c6d6",
   485 => x"feeec600",
   486 => x"c3663c18",
   487 => x"3c66c300",
   488 => x"c3663c18",
   489 => x"18181800",
   490 => x"fe0c1830",
   491 => x"60c0fe00",
   492 => x"3c303030",
   493 => x"30303c00",
   494 => x"c0603018",
   495 => x"0c060300",
   496 => x"3c0c0c0c",
   497 => x"0c0c3c00",
   498 => x"10386cc6",
   499 => x"00000000",
   500 => x"00000000",
   501 => x"000000fe",
   502 => x"18180c00",
   503 => x"00000000",
   504 => x"00003c06",
   505 => x"3e663e00",
   506 => x"60607c66",
   507 => x"66667c00",
   508 => x"00003c60",
   509 => x"60603c00",
   510 => x"06063e66",
   511 => x"66663e00",
   512 => x"00003c66",
   513 => x"7e603c00",
   514 => x"1c307c30",
   515 => x"30303000",
   516 => x"00003e66",
   517 => x"663e063c",
   518 => x"60607c66",
   519 => x"66666600",
   520 => x"18001818",
   521 => x"18180c00",
   522 => x"0c000c0c",
   523 => x"0c0c0c78",
   524 => x"6060666c",
   525 => x"786c6600",
   526 => x"18181818",
   527 => x"18180c00",
   528 => x"0000ecfe",
   529 => x"d6c6c600",
   530 => x"00007c66",
   531 => x"66666600",
   532 => x"00003c66",
   533 => x"66663c00",
   534 => x"00007c66",
   535 => x"667c6060",
   536 => x"00003e66",
   537 => x"663e0606",
   538 => x"00007c66",
   539 => x"60606000",
   540 => x"00003c60",
   541 => x"3c067c00",
   542 => x"30307c30",
   543 => x"30301c00",
   544 => x"00006666",
   545 => x"66663e00",
   546 => x"00006666",
   547 => x"663c1800",
   548 => x"0000c6c6",
   549 => x"d6fe6c00",
   550 => x"0000c66c",
   551 => x"386cc600",
   552 => x"00006666",
   553 => x"663c1830",
   554 => x"00007e0c",
   555 => x"18307e00",
   556 => x"0e181870",
   557 => x"18180e00",
   558 => x"18181818",
   559 => x"18181800",
   560 => x"7018180e",
   561 => x"18187000",
   562 => x"729c0000",
   563 => x"00000000",
   564 => x"fefefefe",
   565 => x"fefefe00",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
   785 => x"00000000",
   786 => x"00000000",
   787 => x"00000000",
   788 => x"00000000",
   789 => x"00000000",
   790 => x"00000000",
   791 => x"00000000",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
   799 => x"00000000",
   800 => x"00000000",
   801 => x"00000000",
   802 => x"00000000",
   803 => x"00000000",
   804 => x"00000000",
   805 => x"00000000",
   806 => x"00000000",
   807 => x"00000000",
   808 => x"00000000",
   809 => x"00000000",
   810 => x"00000000",
   811 => x"00000000",
   812 => x"00000000",
   813 => x"00000000",
   814 => x"00000000",
   815 => x"00000000",
   816 => x"00000000",
   817 => x"00000000",
   818 => x"00000000",
   819 => x"00000000",
   820 => x"00000000",
   821 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

