-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08080f4",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"88907383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02fc050d",
    30 => x"830b85ff",
    31 => x"c48134fc",
    32 => x"0b85ffc0",
    33 => x"8134a080",
    34 => x"81ce2da0",
    35 => x"8083de2d",
    36 => x"80c851a0",
    37 => x"8084922d",
    38 => x"80e551a0",
    39 => x"8084922d",
    40 => x"80ec51a0",
    41 => x"8084922d",
    42 => x"80ec51a0",
    43 => x"8084922d",
    44 => x"80ef51a0",
    45 => x"8084922d",
    46 => x"8a51a080",
    47 => x"84922da0",
    48 => x"8088a051",
    49 => x"a08085f9",
    50 => x"2da08081",
    51 => x"c90402f4",
    52 => x"050dfea0",
    53 => x"800b86ff",
    54 => x"e2802380",
    55 => x"0b86ffe2",
    56 => x"8223800b",
    57 => x"86ffe284",
    58 => x"23800b86",
    59 => x"ffe28823",
    60 => x"800b86ff",
    61 => x"e28a2390",
    62 => x"705353a0",
    63 => x"bf518072",
    64 => x"70840554",
    65 => x"0cff1151",
    66 => x"708025f2",
    67 => x"38bc0b86",
    68 => x"ffe19223",
    69 => x"81d40b86",
    70 => x"ffe19423",
    71 => x"80d9810b",
    72 => x"86ffe18e",
    73 => x"23e9c10b",
    74 => x"86ffe190",
    75 => x"2386ff0b",
    76 => x"86ffe380",
    77 => x"239fff0b",
    78 => x"86ffe382",
    79 => x"2381e00b",
    80 => x"84889023",
    81 => x"900b902c",
    82 => x"51708488",
    83 => x"922381e2",
    84 => x"0b848894",
    85 => x"23728488",
    86 => x"9623ff0b",
    87 => x"84889823",
    88 => x"fe0b8488",
    89 => x"9a238488",
    90 => x"900b902c",
    91 => x"527186ff",
    92 => x"e1802384",
    93 => x"88905170",
    94 => x"86ffe182",
    95 => x"23800b86",
    96 => x"ffe18823",
    97 => x"fe87900b",
    98 => x"86ffe196",
    99 => x"23800b84",
   100 => x"88a00c80",
   101 => x"0b8488a4",
   102 => x"0c028c05",
   103 => x"0d0402f8",
   104 => x"050d8488",
   105 => x"a4081010",
   106 => x"8488a408",
   107 => x"05709029",
   108 => x"8488a008",
   109 => x"0584c011",
   110 => x"51525280",
   111 => x"52717134",
   112 => x"71811234",
   113 => x"71821234",
   114 => x"71831234",
   115 => x"80d01181",
   116 => x"13535181",
   117 => x"ff7225e5",
   118 => x"38028805",
   119 => x"0d0402f4",
   120 => x"050d9053",
   121 => x"a0bf5272",
   122 => x"84147108",
   123 => x"8105720c",
   124 => x"ff145454",
   125 => x"51807224",
   126 => x"e9387284",
   127 => x"14710881",
   128 => x"05720cff",
   129 => x"14545451",
   130 => x"718025db",
   131 => x"38a08083",
   132 => x"e20402e8",
   133 => x"050d7756",
   134 => x"9f762581",
   135 => x"8d388488",
   136 => x"a4087010",
   137 => x"10117081",
   138 => x"80298488",
   139 => x"a0080584",
   140 => x"c0117910",
   141 => x"1010a080",
   142 => x"86b00570",
   143 => x"70840552",
   144 => x"08710852",
   145 => x"54555154",
   146 => x"55557072",
   147 => x"3470882c",
   148 => x"5372ffb0",
   149 => x"13347090",
   150 => x"2c5372fe",
   151 => x"e0133470",
   152 => x"982c5170",
   153 => x"fe901334",
   154 => x"73fdc013",
   155 => x"3473882c",
   156 => x"5372fcf0",
   157 => x"13347390",
   158 => x"2c5170fc",
   159 => x"a0133473",
   160 => x"982c5473",
   161 => x"fbd01334",
   162 => x"758a2eab",
   163 => x"388488a0",
   164 => x"08810584",
   165 => x"88a00c84",
   166 => x"88a00880",
   167 => x"d02e9838",
   168 => x"74992eac",
   169 => x"38029805",
   170 => x"0d048488",
   171 => x"a4085575",
   172 => x"8a2e0981",
   173 => x"06d73881",
   174 => x"158488a4",
   175 => x"0c800b84",
   176 => x"88a00c84",
   177 => x"88a40855",
   178 => x"74992e09",
   179 => x"8106d638",
   180 => x"900b9480",
   181 => x"1154529f",
   182 => x"9f517270",
   183 => x"84055408",
   184 => x"72708405",
   185 => x"540cff11",
   186 => x"51708025",
   187 => x"ed38980b",
   188 => x"8488a40c",
   189 => x"0298050d",
   190 => x"0402dc05",
   191 => x"0d7a5877",
   192 => x"70840559",
   193 => x"08578059",
   194 => x"76982a77",
   195 => x"882b5856",
   196 => x"75802e81",
   197 => x"9b389f76",
   198 => x"25819a38",
   199 => x"8488a408",
   200 => x"70101011",
   201 => x"70818029",
   202 => x"8488a008",
   203 => x"0584c011",
   204 => x"79101010",
   205 => x"a08086b0",
   206 => x"05707084",
   207 => x"05520871",
   208 => x"08525455",
   209 => x"51545555",
   210 => x"70723470",
   211 => x"882c5372",
   212 => x"ffb01334",
   213 => x"70902c53",
   214 => x"72fee013",
   215 => x"3470982c",
   216 => x"5170fe90",
   217 => x"133473fd",
   218 => x"c0133473",
   219 => x"882c5372",
   220 => x"fcf01334",
   221 => x"73902c51",
   222 => x"70fca013",
   223 => x"3473982c",
   224 => x"5473fbd0",
   225 => x"1334758a",
   226 => x"2eb83884",
   227 => x"88a00881",
   228 => x"058488a0",
   229 => x"0c8488a0",
   230 => x"0880d02e",
   231 => x"a5387499",
   232 => x"2eb93881",
   233 => x"19598379",
   234 => x"25fedd38",
   235 => x"75fed038",
   236 => x"02a4050d",
   237 => x"048488a4",
   238 => x"0855758a",
   239 => x"2e098106",
   240 => x"ca388115",
   241 => x"8488a40c",
   242 => x"800b8488",
   243 => x"a00c8488",
   244 => x"a4085574",
   245 => x"992e0981",
   246 => x"06c93890",
   247 => x"0b948011",
   248 => x"54529f9f",
   249 => x"51727084",
   250 => x"05540872",
   251 => x"70840554",
   252 => x"0cff1151",
   253 => x"708025ed",
   254 => x"38980b84",
   255 => x"88a40c81",
   256 => x"19598379",
   257 => x"25fe8138",
   258 => x"a08087ac",
   259 => x"04000000",
   260 => x"00ffffff",
   261 => x"ff00ffff",
   262 => x"ffff00ff",
   263 => x"ffffff00",
   264 => x"48656c6c",
   265 => x"6f2c2077",
   266 => x"6f726c64",
   267 => x"210a0000",
   268 => x"00000000",
   269 => x"00000000",
   270 => x"18181818",
   271 => x"18001800",
   272 => x"6c6c0000",
   273 => x"00000000",
   274 => x"6c6cfe6c",
   275 => x"fe6c6c00",
   276 => x"183e603c",
   277 => x"067c1800",
   278 => x"0066acd8",
   279 => x"366acc00",
   280 => x"386c6876",
   281 => x"dcce7b00",
   282 => x"18183000",
   283 => x"00000000",
   284 => x"0c183030",
   285 => x"30180c00",
   286 => x"30180c0c",
   287 => x"0c183000",
   288 => x"00663cff",
   289 => x"3c660000",
   290 => x"0018187e",
   291 => x"18180000",
   292 => x"00000000",
   293 => x"00181830",
   294 => x"0000007e",
   295 => x"00000000",
   296 => x"00000000",
   297 => x"00181800",
   298 => x"03060c18",
   299 => x"3060c000",
   300 => x"3c666e7e",
   301 => x"76663c00",
   302 => x"18387818",
   303 => x"18181800",
   304 => x"3c66060c",
   305 => x"18307e00",
   306 => x"3c66061c",
   307 => x"06663c00",
   308 => x"1c3c6ccc",
   309 => x"fe0c0c00",
   310 => x"7e607c06",
   311 => x"06663c00",
   312 => x"1c30607c",
   313 => x"66663c00",
   314 => x"7e06060c",
   315 => x"18181800",
   316 => x"3c66663c",
   317 => x"66663c00",
   318 => x"3c66663e",
   319 => x"060c3800",
   320 => x"00181800",
   321 => x"00181800",
   322 => x"00181800",
   323 => x"00181830",
   324 => x"00061860",
   325 => x"18060000",
   326 => x"00007e00",
   327 => x"7e000000",
   328 => x"00601806",
   329 => x"18600000",
   330 => x"3c66060c",
   331 => x"18001800",
   332 => x"7cc6ded6",
   333 => x"dec07800",
   334 => x"3c66667e",
   335 => x"66666600",
   336 => x"7c66667c",
   337 => x"66667c00",
   338 => x"1e306060",
   339 => x"60301e00",
   340 => x"786c6666",
   341 => x"666c7800",
   342 => x"7e606078",
   343 => x"60607e00",
   344 => x"7e606078",
   345 => x"60606000",
   346 => x"3c66606e",
   347 => x"66663e00",
   348 => x"6666667e",
   349 => x"66666600",
   350 => x"3c181818",
   351 => x"18183c00",
   352 => x"06060606",
   353 => x"06663c00",
   354 => x"c6ccd8f0",
   355 => x"d8ccc600",
   356 => x"60606060",
   357 => x"60607e00",
   358 => x"c6eefed6",
   359 => x"c6c6c600",
   360 => x"c6e6f6de",
   361 => x"cec6c600",
   362 => x"3c666666",
   363 => x"66663c00",
   364 => x"7c66667c",
   365 => x"60606000",
   366 => x"78cccccc",
   367 => x"ccdc7e00",
   368 => x"7c66667c",
   369 => x"6c666600",
   370 => x"3c66703c",
   371 => x"0e663c00",
   372 => x"7e181818",
   373 => x"18181800",
   374 => x"66666666",
   375 => x"66663c00",
   376 => x"66666666",
   377 => x"3c3c1800",
   378 => x"c6c6c6d6",
   379 => x"feeec600",
   380 => x"c3663c18",
   381 => x"3c66c300",
   382 => x"c3663c18",
   383 => x"18181800",
   384 => x"fe0c1830",
   385 => x"60c0fe00",
   386 => x"3c303030",
   387 => x"30303c00",
   388 => x"c0603018",
   389 => x"0c060300",
   390 => x"3c0c0c0c",
   391 => x"0c0c3c00",
   392 => x"10386cc6",
   393 => x"00000000",
   394 => x"00000000",
   395 => x"000000fe",
   396 => x"18180c00",
   397 => x"00000000",
   398 => x"00003c06",
   399 => x"3e663e00",
   400 => x"60607c66",
   401 => x"66667c00",
   402 => x"00003c60",
   403 => x"60603c00",
   404 => x"06063e66",
   405 => x"66663e00",
   406 => x"00003c66",
   407 => x"7e603c00",
   408 => x"1c307c30",
   409 => x"30303000",
   410 => x"00003e66",
   411 => x"663e063c",
   412 => x"60607c66",
   413 => x"66666600",
   414 => x"18001818",
   415 => x"18180c00",
   416 => x"0c000c0c",
   417 => x"0c0c0c78",
   418 => x"6060666c",
   419 => x"786c6600",
   420 => x"18181818",
   421 => x"18180c00",
   422 => x"0000ecfe",
   423 => x"d6c6c600",
   424 => x"00007c66",
   425 => x"66666600",
   426 => x"00003c66",
   427 => x"66663c00",
   428 => x"00007c66",
   429 => x"667c6060",
   430 => x"00003e66",
   431 => x"663e0606",
   432 => x"00007c66",
   433 => x"60606000",
   434 => x"00003c60",
   435 => x"3c067c00",
   436 => x"30307c30",
   437 => x"30301c00",
   438 => x"00006666",
   439 => x"66663e00",
   440 => x"00006666",
   441 => x"663c1800",
   442 => x"0000c6c6",
   443 => x"d6fe6c00",
   444 => x"0000c66c",
   445 => x"386cc600",
   446 => x"00006666",
   447 => x"663c1830",
   448 => x"00007e0c",
   449 => x"18307e00",
   450 => x"0e181870",
   451 => x"18180e00",
   452 => x"18181818",
   453 => x"18181800",
   454 => x"7018180e",
   455 => x"18187000",
   456 => x"729c0000",
   457 => x"00000000",
   458 => x"fefefefe",
   459 => x"fefefe00",
   460 => x"00000000",
   461 => x"00000000",
   462 => x"00000000",
   463 => x"00000000",
   464 => x"00000000",
   465 => x"00000000",
   466 => x"00000000",
   467 => x"00000000",
   468 => x"00000000",
   469 => x"00000000",
   470 => x"00000000",
   471 => x"00000000",
   472 => x"00000000",
   473 => x"00000000",
   474 => x"00000000",
   475 => x"00000000",
   476 => x"00000000",
   477 => x"00000000",
   478 => x"00000000",
   479 => x"00000000",
   480 => x"00000000",
   481 => x"00000000",
   482 => x"00000000",
   483 => x"00000000",
   484 => x"00000000",
   485 => x"00000000",
   486 => x"00000000",
   487 => x"00000000",
   488 => x"00000000",
   489 => x"00000000",
   490 => x"00000000",
   491 => x"00000000",
   492 => x"00000000",
   493 => x"00000000",
   494 => x"00000000",
   495 => x"00000000",
   496 => x"00000000",
   497 => x"00000000",
   498 => x"00000000",
   499 => x"00000000",
   500 => x"00000000",
   501 => x"00000000",
   502 => x"00000000",
   503 => x"00000000",
   504 => x"00000000",
   505 => x"00000000",
   506 => x"00000000",
   507 => x"00000000",
   508 => x"00000000",
   509 => x"00000000",
   510 => x"00000000",
   511 => x"00000000",
   512 => x"00000000",
   513 => x"00000000",
   514 => x"00000000",
   515 => x"00000000",
   516 => x"00000000",
   517 => x"00000000",
   518 => x"00000000",
   519 => x"00000000",
   520 => x"00000000",
   521 => x"00000000",
   522 => x"00000000",
   523 => x"00000000",
   524 => x"00000000",
   525 => x"00000000",
   526 => x"00000000",
   527 => x"00000000",
   528 => x"00000000",
   529 => x"00000000",
   530 => x"00000000",
   531 => x"00000000",
   532 => x"00000000",
   533 => x"00000000",
   534 => x"00000000",
   535 => x"00000000",
   536 => x"00000000",
   537 => x"00000000",
   538 => x"00000000",
   539 => x"00000000",
   540 => x"00000000",
   541 => x"00000000",
   542 => x"00000000",
   543 => x"00000000",
   544 => x"00000000",
   545 => x"00000000",
   546 => x"00000000",
   547 => x"00000000",
   548 => x"00000000",
   549 => x"00000000",
   550 => x"00000000",
   551 => x"00000000",
   552 => x"00000000",
   553 => x"00000000",
   554 => x"00000000",
   555 => x"00000000",
   556 => x"00000000",
   557 => x"00000000",
   558 => x"00000000",
   559 => x"00000000",
   560 => x"00000000",
   561 => x"00000000",
   562 => x"00000000",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

