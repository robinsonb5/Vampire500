-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08094e5",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"95f07383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02f8050d",
    30 => x"028f05a0",
    31 => x"8080b42d",
    32 => x"52ff8408",
    33 => x"70882a70",
    34 => x"81065151",
    35 => x"5170802e",
    36 => x"f03871ff",
    37 => x"840c0288",
    38 => x"050d0402",
    39 => x"f4050d74",
    40 => x"5372a080",
    41 => x"80b42d70",
    42 => x"81ff0652",
    43 => x"5270802e",
    44 => x"a3387181",
    45 => x"ff068114",
    46 => x"5452ff84",
    47 => x"0870882a",
    48 => x"70810651",
    49 => x"51517080",
    50 => x"2ef03871",
    51 => x"ff840ca0",
    52 => x"8081a104",
    53 => x"028c050d",
    54 => x"0402f805",
    55 => x"0d028f05",
    56 => x"a08080b4",
    57 => x"2d52ff84",
    58 => x"0870882a",
    59 => x"70810651",
    60 => x"51517080",
    61 => x"2ef03871",
    62 => x"ff840c02",
    63 => x"88050d04",
    64 => x"02d0050d",
    65 => x"02b405a0",
    66 => x"8081d971",
    67 => x"70840553",
    68 => x"085c5c58",
    69 => x"807a7081",
    70 => x"055ca080",
    71 => x"80b42d54",
    72 => x"5972792e",
    73 => x"82cc3872",
    74 => x"a52e0981",
    75 => x"0682ab38",
    76 => x"79708105",
    77 => x"5ba08080",
    78 => x"b42d5372",
    79 => x"80e42e9f",
    80 => x"387280e4",
    81 => x"248d3872",
    82 => x"80e32e81",
    83 => x"c438a080",
    84 => x"84a30472",
    85 => x"80f32e81",
    86 => x"8d38a080",
    87 => x"84a30477",
    88 => x"84197108",
    89 => x"a0809ee0",
    90 => x"0ba0809e",
    91 => x"90595a56",
    92 => x"59538056",
    93 => x"73762e09",
    94 => x"81069538",
    95 => x"b00ba080",
    96 => x"9e900ba0",
    97 => x"8080c92d",
    98 => x"811555a0",
    99 => x"8083b804",
   100 => x"738f06a0",
   101 => x"80968005",
   102 => x"5372a080",
   103 => x"80b42d75",
   104 => x"70810557",
   105 => x"a08080c9",
   106 => x"2d73842a",
   107 => x"5473e138",
   108 => x"74a0809e",
   109 => x"902e9c38",
   110 => x"ff155574",
   111 => x"a08080b4",
   112 => x"2d777081",
   113 => x"0559a080",
   114 => x"80c92d81",
   115 => x"1656a080",
   116 => x"83b00480",
   117 => x"77a08080",
   118 => x"c92d75a0",
   119 => x"809ee056",
   120 => x"54a08084",
   121 => x"b7047784",
   122 => x"19710857",
   123 => x"59538075",
   124 => x"a08080b4",
   125 => x"2d545472",
   126 => x"742ebc38",
   127 => x"81147016",
   128 => x"70a08080",
   129 => x"b42d5154",
   130 => x"5472f138",
   131 => x"a08084b7",
   132 => x"04778419",
   133 => x"8312a080",
   134 => x"80b42d52",
   135 => x"5953a080",
   136 => x"84da0480",
   137 => x"52a5517a",
   138 => x"2d805272",
   139 => x"517a2d82",
   140 => x"1959a080",
   141 => x"84e30473",
   142 => x"ff155553",
   143 => x"807325a3",
   144 => x"38747081",
   145 => x"0556a080",
   146 => x"80b42d53",
   147 => x"80527251",
   148 => x"7a2d8119",
   149 => x"59a08084",
   150 => x"b7048052",
   151 => x"72517a2d",
   152 => x"81195979",
   153 => x"7081055b",
   154 => x"a08080b4",
   155 => x"2d5372fd",
   156 => x"b63878a0",
   157 => x"809e800c",
   158 => x"02b0050d",
   159 => x"0402f405",
   160 => x"0d747671",
   161 => x"81ff06c8",
   162 => x"0c5353a0",
   163 => x"809fa008",
   164 => x"85387189",
   165 => x"2b527198",
   166 => x"2ac80c71",
   167 => x"902a7081",
   168 => x"ff06c80c",
   169 => x"5171882a",
   170 => x"7081ff06",
   171 => x"c80c5171",
   172 => x"81ff06c8",
   173 => x"0c72902a",
   174 => x"7081ff06",
   175 => x"c80c51c8",
   176 => x"087081ff",
   177 => x"06515182",
   178 => x"b8bf5270",
   179 => x"81ff2e09",
   180 => x"81069438",
   181 => x"81ff0bc8",
   182 => x"0cc80870",
   183 => x"81ff06ff",
   184 => x"14545151",
   185 => x"71e53870",
   186 => x"a0809e80",
   187 => x"0c028c05",
   188 => x"0d0402fc",
   189 => x"050d81c7",
   190 => x"5181ff0b",
   191 => x"c80cff11",
   192 => x"51708025",
   193 => x"f4380284",
   194 => x"050d0402",
   195 => x"f0050da0",
   196 => x"8085f22d",
   197 => x"819c9f53",
   198 => x"805287fc",
   199 => x"80f751a0",
   200 => x"8084fd2d",
   201 => x"a0809e80",
   202 => x"0854a080",
   203 => x"9e800881",
   204 => x"2e098106",
   205 => x"ab3881ff",
   206 => x"0bc80c82",
   207 => x"0a52849c",
   208 => x"80e951a0",
   209 => x"8084fd2d",
   210 => x"a0809e80",
   211 => x"088d3881",
   212 => x"ff0bc80c",
   213 => x"7353a080",
   214 => x"86e704a0",
   215 => x"8085f22d",
   216 => x"ff135372",
   217 => x"ffb23872",
   218 => x"a0809e80",
   219 => x"0c029005",
   220 => x"0d0402f4",
   221 => x"050d81ff",
   222 => x"0bc80c93",
   223 => x"53805287",
   224 => x"fc80c151",
   225 => x"a08084fd",
   226 => x"2da0809e",
   227 => x"80088d38",
   228 => x"81ff0bc8",
   229 => x"0c8153a0",
   230 => x"8087a704",
   231 => x"a08085f2",
   232 => x"2dff1353",
   233 => x"72d73872",
   234 => x"a0809e80",
   235 => x"0c028c05",
   236 => x"0d0402f0",
   237 => x"050da080",
   238 => x"85f22d83",
   239 => x"aa52849c",
   240 => x"80c851a0",
   241 => x"8084fd2d",
   242 => x"a0809e80",
   243 => x"08812e09",
   244 => x"81068e38",
   245 => x"cc0883ff",
   246 => x"ff065372",
   247 => x"83aa2ea3",
   248 => x"38a08086",
   249 => x"f22da080",
   250 => x"87fc0481",
   251 => x"54a08089",
   252 => x"9304a080",
   253 => x"969451a0",
   254 => x"8082802d",
   255 => x"8054a080",
   256 => x"89930481",
   257 => x"ff0bc80c",
   258 => x"b153a080",
   259 => x"868b2da0",
   260 => x"809e8008",
   261 => x"802e80e2",
   262 => x"38805287",
   263 => x"fc80fa51",
   264 => x"a08084fd",
   265 => x"2da0809e",
   266 => x"8008bf38",
   267 => x"a0809e80",
   268 => x"0852a080",
   269 => x"96b051a0",
   270 => x"8082802d",
   271 => x"81ff0bc8",
   272 => x"0cc80881",
   273 => x"ff067053",
   274 => x"a08096bc",
   275 => x"5254a080",
   276 => x"82802dcc",
   277 => x"0874862a",
   278 => x"70810670",
   279 => x"57515153",
   280 => x"72802eaf",
   281 => x"38a08087",
   282 => x"eb04a080",
   283 => x"9e800852",
   284 => x"a08096b0",
   285 => x"51a08082",
   286 => x"802d7282",
   287 => x"2efef338",
   288 => x"ff135372",
   289 => x"ff8438a0",
   290 => x"8096cc51",
   291 => x"a080819b",
   292 => x"2d725473",
   293 => x"a0809e80",
   294 => x"0c029005",
   295 => x"0d0402f4",
   296 => x"050d810b",
   297 => x"a0809fa0",
   298 => x"0cc40870",
   299 => x"8f2a7081",
   300 => x"06515153",
   301 => x"72f33872",
   302 => x"c40ca080",
   303 => x"85f22dc4",
   304 => x"08708f2a",
   305 => x"70810651",
   306 => x"515372f3",
   307 => x"38810bc4",
   308 => x"0c875380",
   309 => x"5284d480",
   310 => x"c051a080",
   311 => x"84fd2da0",
   312 => x"809e8008",
   313 => x"812e0981",
   314 => x"068738a0",
   315 => x"809e8008",
   316 => x"53a08096",
   317 => x"e451a080",
   318 => x"819b2d72",
   319 => x"822e0981",
   320 => x"069238a0",
   321 => x"8096f851",
   322 => x"a080819b",
   323 => x"2d8053a0",
   324 => x"808b8404",
   325 => x"ff135372",
   326 => x"ffb938a0",
   327 => x"80979851",
   328 => x"a080819b",
   329 => x"2da08087",
   330 => x"b22da080",
   331 => x"9e8008a0",
   332 => x"809fa00c",
   333 => x"a0809e80",
   334 => x"08802e8b",
   335 => x"38a08097",
   336 => x"b451a080",
   337 => x"819b2da0",
   338 => x"8097c851",
   339 => x"a080819b",
   340 => x"2d815287",
   341 => x"fc80d051",
   342 => x"a08084fd",
   343 => x"2d81ff0b",
   344 => x"c80cc408",
   345 => x"708f2a70",
   346 => x"81065151",
   347 => x"5372f338",
   348 => x"72c40c81",
   349 => x"ff0bc80c",
   350 => x"a08097d8",
   351 => x"51a08081",
   352 => x"9b2d8153",
   353 => x"72a0809e",
   354 => x"800c028c",
   355 => x"050d0480",
   356 => x"0ba0809e",
   357 => x"800c0402",
   358 => x"e0050d79",
   359 => x"7b575780",
   360 => x"58c40870",
   361 => x"8f2a7081",
   362 => x"06515154",
   363 => x"73f33882",
   364 => x"810bc40c",
   365 => x"81ff0bc8",
   366 => x"0c765287",
   367 => x"fc80d151",
   368 => x"a08084fd",
   369 => x"2d80dbc6",
   370 => x"df55a080",
   371 => x"9e800880",
   372 => x"2e9838a0",
   373 => x"809e8008",
   374 => x"537652a0",
   375 => x"8097e451",
   376 => x"a0808280",
   377 => x"2da0808c",
   378 => x"b60481ff",
   379 => x"0bc80cc8",
   380 => x"087081ff",
   381 => x"06515473",
   382 => x"81fe2e09",
   383 => x"81069b38",
   384 => x"80ff55cc",
   385 => x"08767084",
   386 => x"05580cff",
   387 => x"15557480",
   388 => x"25f13881",
   389 => x"58a0808c",
   390 => x"a004ff15",
   391 => x"5574cb38",
   392 => x"81ff0bc8",
   393 => x"0cc40870",
   394 => x"8f2a7081",
   395 => x"06515154",
   396 => x"73f33873",
   397 => x"c40c77a0",
   398 => x"809e800c",
   399 => x"02a0050d",
   400 => x"0402f405",
   401 => x"0d747088",
   402 => x"2a83fe80",
   403 => x"06707298",
   404 => x"2a077288",
   405 => x"2b87fc80",
   406 => x"80067398",
   407 => x"2b81f00a",
   408 => x"06717307",
   409 => x"07a0809e",
   410 => x"800c5651",
   411 => x"5351028c",
   412 => x"050d0402",
   413 => x"f4050d02",
   414 => x"92052270",
   415 => x"882a7188",
   416 => x"2b077083",
   417 => x"ffff06a0",
   418 => x"809e800c",
   419 => x"5252028c",
   420 => x"050d0402",
   421 => x"f8050d73",
   422 => x"70902b71",
   423 => x"902a07a0",
   424 => x"809e800c",
   425 => x"52028805",
   426 => x"0d0402f4",
   427 => x"050d7476",
   428 => x"52538071",
   429 => x"25903870",
   430 => x"52727084",
   431 => x"055408ff",
   432 => x"13535171",
   433 => x"f438028c",
   434 => x"050d0402",
   435 => x"d8050d7b",
   436 => x"7d5b5681",
   437 => x"0ba08098",
   438 => x"84595783",
   439 => x"59770876",
   440 => x"0c750878",
   441 => x"08565473",
   442 => x"752e9238",
   443 => x"75085374",
   444 => x"52a08098",
   445 => x"9451a080",
   446 => x"82802d80",
   447 => x"57795275",
   448 => x"51a0808d",
   449 => x"aa2d7508",
   450 => x"5473752e",
   451 => x"92387508",
   452 => x"537452a0",
   453 => x"8098d451",
   454 => x"a0808280",
   455 => x"2d8057ff",
   456 => x"19841959",
   457 => x"59788025",
   458 => x"ffb33876",
   459 => x"a0809e80",
   460 => x"0c02a805",
   461 => x"0d0402ec",
   462 => x"050d7654",
   463 => x"815585aa",
   464 => x"d5aad574",
   465 => x"0cfad5aa",
   466 => x"d5aa0b8c",
   467 => x"150ccc74",
   468 => x"a08080c9",
   469 => x"2db30b8f",
   470 => x"15a08080",
   471 => x"c92d7308",
   472 => x"5372fce2",
   473 => x"d5aad52e",
   474 => x"90387308",
   475 => x"52a08099",
   476 => x"9451a080",
   477 => x"82802d80",
   478 => x"558c1408",
   479 => x"5372fad5",
   480 => x"aad4b32e",
   481 => x"91388c14",
   482 => x"0852a080",
   483 => x"99d051a0",
   484 => x"8082802d",
   485 => x"80557752",
   486 => x"7351a080",
   487 => x"8daa2d73",
   488 => x"085372fc",
   489 => x"e2d5aad5",
   490 => x"2e903873",
   491 => x"0852a080",
   492 => x"9a8c51a0",
   493 => x"8082802d",
   494 => x"80558c14",
   495 => x"085372fa",
   496 => x"d5aad4b3",
   497 => x"2e91388c",
   498 => x"140852a0",
   499 => x"809ac851",
   500 => x"a0808280",
   501 => x"2d805574",
   502 => x"a0809e80",
   503 => x"0c029405",
   504 => x"0d0402c8",
   505 => x"050d7f5c",
   506 => x"800ba080",
   507 => x"9b84525b",
   508 => x"a0808280",
   509 => x"2d80e1b3",
   510 => x"578e5d76",
   511 => x"598fffff",
   512 => x"5a76bfff",
   513 => x"ff067710",
   514 => x"70962a70",
   515 => x"81065157",
   516 => x"58587480",
   517 => x"2e853876",
   518 => x"81075776",
   519 => x"952a7081",
   520 => x"06515574",
   521 => x"802e8538",
   522 => x"76813257",
   523 => x"76bfffff",
   524 => x"06788429",
   525 => x"1d79710c",
   526 => x"56708429",
   527 => x"1d56750c",
   528 => x"76107096",
   529 => x"2a708106",
   530 => x"51565774",
   531 => x"802e8538",
   532 => x"76810757",
   533 => x"76952a70",
   534 => x"81065155",
   535 => x"74802e85",
   536 => x"38768132",
   537 => x"57ff1a5a",
   538 => x"798025ff",
   539 => x"94387857",
   540 => x"8fffff5a",
   541 => x"76bfffff",
   542 => x"06771070",
   543 => x"962a7081",
   544 => x"06515758",
   545 => x"5674802e",
   546 => x"85387681",
   547 => x"07577695",
   548 => x"2a708106",
   549 => x"51557480",
   550 => x"2e853876",
   551 => x"81325776",
   552 => x"bfffff06",
   553 => x"7684291d",
   554 => x"7008575a",
   555 => x"5874762e",
   556 => x"a738807b",
   557 => x"53a0809b",
   558 => x"98525ea0",
   559 => x"8082802d",
   560 => x"78085475",
   561 => x"537552a0",
   562 => x"809bac51",
   563 => x"a0808280",
   564 => x"2d7d5ba0",
   565 => x"8091db04",
   566 => x"811b5b77",
   567 => x"84291c70",
   568 => x"08565674",
   569 => x"782ea738",
   570 => x"807b53a0",
   571 => x"809b9852",
   572 => x"5ea08082",
   573 => x"802d7508",
   574 => x"54775377",
   575 => x"52a0809b",
   576 => x"ac51a080",
   577 => x"82802d7d",
   578 => x"5ba08092",
   579 => x"9104811b",
   580 => x"5b761070",
   581 => x"962a7081",
   582 => x"06515657",
   583 => x"74802e85",
   584 => x"38768107",
   585 => x"5776952a",
   586 => x"70810651",
   587 => x"5574802e",
   588 => x"85387681",
   589 => x"3257ff1a",
   590 => x"5a798025",
   591 => x"feb638ff",
   592 => x"1d5d7cfd",
   593 => x"b6387da0",
   594 => x"809e800c",
   595 => x"02b8050d",
   596 => x"0402cc05",
   597 => x"0d7e5c81",
   598 => x"5b805a80",
   599 => x"c07b585d",
   600 => x"85ada989",
   601 => x"bb7c0c7a",
   602 => x"56815897",
   603 => x"55767807",
   604 => x"822b7c11",
   605 => x"515485ad",
   606 => x"a989bb74",
   607 => x"0c7710ff",
   608 => x"16565874",
   609 => x"8025e638",
   610 => x"76108117",
   611 => x"57579876",
   612 => x"25d7387f",
   613 => x"527b51a0",
   614 => x"808daa2d",
   615 => x"8157ff87",
   616 => x"87a5c37c",
   617 => x"0c975680",
   618 => x"77822b7d",
   619 => x"11700857",
   620 => x"575a5873",
   621 => x"ff8787a5",
   622 => x"c32e0981",
   623 => x"068a3879",
   624 => x"77075aa0",
   625 => x"8093e504",
   626 => x"74085473",
   627 => x"85ada989",
   628 => x"bb2e9238",
   629 => x"77750854",
   630 => x"7953a080",
   631 => x"9bd4525b",
   632 => x"a0808280",
   633 => x"2d7610ff",
   634 => x"17575775",
   635 => x"8025ffb7",
   636 => x"3879802e",
   637 => x"ba387982",
   638 => x"2b52a080",
   639 => x"9bf451a0",
   640 => x"8082802d",
   641 => x"79992a81",
   642 => x"32708106",
   643 => x"70098105",
   644 => x"70720770",
   645 => x"09709f2c",
   646 => x"60067f10",
   647 => x"87fffffe",
   648 => x"0663812c",
   649 => x"44404051",
   650 => x"51565155",
   651 => x"79d6387a",
   652 => x"09810570",
   653 => x"7c079f2a",
   654 => x"51547cbf",
   655 => x"24903873",
   656 => x"802e8b38",
   657 => x"a0809c8c",
   658 => x"51a08082",
   659 => x"802d7c52",
   660 => x"a0809cd8",
   661 => x"51a08082",
   662 => x"802d7aa0",
   663 => x"809e800c",
   664 => x"02b4050d",
   665 => x"0402f805",
   666 => x"0d88bd0b",
   667 => x"ff880ca0",
   668 => x"80528051",
   669 => x"a0808dcb",
   670 => x"2da0809e",
   671 => x"8008802e",
   672 => x"8b38a080",
   673 => x"9d9451a0",
   674 => x"8082802d",
   675 => x"a0805280",
   676 => x"51a0808e",
   677 => x"b62da080",
   678 => x"9e800880",
   679 => x"2e8b38a0",
   680 => x"809db851",
   681 => x"a0808280",
   682 => x"2da08052",
   683 => x"8051a080",
   684 => x"92d12da0",
   685 => x"809e8008",
   686 => x"802e8b38",
   687 => x"a0809dd4",
   688 => x"51a08082",
   689 => x"802d8051",
   690 => x"a0808fe2",
   691 => x"2da0809e",
   692 => x"8008802e",
   693 => x"8b38a080",
   694 => x"9dec51a0",
   695 => x"8082802d",
   696 => x"a08099cc",
   697 => x"51a08082",
   698 => x"802da080",
   699 => x"94ef0400",
   700 => x"00ffffff",
   701 => x"ff00ffff",
   702 => x"ffff00ff",
   703 => x"ffffff00",
   704 => x"30313233",
   705 => x"34353637",
   706 => x"38394142",
   707 => x"43444546",
   708 => x"00000000",
   709 => x"53444843",
   710 => x"20496e69",
   711 => x"7469616c",
   712 => x"697a6174",
   713 => x"696f6e20",
   714 => x"6572726f",
   715 => x"72210a00",
   716 => x"434d4435",
   717 => x"38202564",
   718 => x"0a202000",
   719 => x"434d4435",
   720 => x"385f3220",
   721 => x"25640a20",
   722 => x"20000000",
   723 => x"44657465",
   724 => x"726d696e",
   725 => x"65642053",
   726 => x"44484320",
   727 => x"73746174",
   728 => x"75730a00",
   729 => x"53656e74",
   730 => x"20726573",
   731 => x"65742063",
   732 => x"6f6d6d61",
   733 => x"6e640a00",
   734 => x"53442063",
   735 => x"61726420",
   736 => x"696e6974",
   737 => x"69616c69",
   738 => x"7a617469",
   739 => x"6f6e2065",
   740 => x"72726f72",
   741 => x"210a0000",
   742 => x"43617264",
   743 => x"20726573",
   744 => x"706f6e64",
   745 => x"65642074",
   746 => x"6f207265",
   747 => x"7365740a",
   748 => x"00000000",
   749 => x"53444843",
   750 => x"20636172",
   751 => x"64206465",
   752 => x"74656374",
   753 => x"65640a00",
   754 => x"53656e64",
   755 => x"696e6720",
   756 => x"636d6431",
   757 => x"360a0000",
   758 => x"496e6974",
   759 => x"20646f6e",
   760 => x"650a0000",
   761 => x"52656164",
   762 => x"20636f6d",
   763 => x"6d616e64",
   764 => x"20666169",
   765 => x"6c656420",
   766 => x"61742025",
   767 => x"64202825",
   768 => x"64290a00",
   769 => x"00000000",
   770 => x"55555555",
   771 => x"aaaaaaaa",
   772 => x"ffffffff",
   773 => x"53616e69",
   774 => x"74792063",
   775 => x"6865636b",
   776 => x"20666169",
   777 => x"6c656420",
   778 => x"28626566",
   779 => x"6f726520",
   780 => x"63616368",
   781 => x"65207265",
   782 => x"66726573",
   783 => x"6829206f",
   784 => x"6e203078",
   785 => x"25642028",
   786 => x"676f7420",
   787 => x"30782564",
   788 => x"290a0000",
   789 => x"53616e69",
   790 => x"74792063",
   791 => x"6865636b",
   792 => x"20666169",
   793 => x"6c656420",
   794 => x"28616674",
   795 => x"65722063",
   796 => x"61636865",
   797 => x"20726566",
   798 => x"72657368",
   799 => x"29206f6e",
   800 => x"20307825",
   801 => x"64202867",
   802 => x"6f742030",
   803 => x"78256429",
   804 => x"0a000000",
   805 => x"42797465",
   806 => x"20636865",
   807 => x"636b2066",
   808 => x"61696c65",
   809 => x"64202862",
   810 => x"65666f72",
   811 => x"65206361",
   812 => x"63686520",
   813 => x"72656672",
   814 => x"65736829",
   815 => x"20617420",
   816 => x"30202867",
   817 => x"6f742030",
   818 => x"78256429",
   819 => x"0a000000",
   820 => x"42797465",
   821 => x"20636865",
   822 => x"636b2066",
   823 => x"61696c65",
   824 => x"64202862",
   825 => x"65666f72",
   826 => x"65206361",
   827 => x"63686520",
   828 => x"72656672",
   829 => x"65736829",
   830 => x"20617420",
   831 => x"33202867",
   832 => x"6f742030",
   833 => x"78256429",
   834 => x"0a000000",
   835 => x"42797465",
   836 => x"20636865",
   837 => x"636b2066",
   838 => x"61696c65",
   839 => x"64202861",
   840 => x"66746572",
   841 => x"20636163",
   842 => x"68652072",
   843 => x"65667265",
   844 => x"73682920",
   845 => x"61742030",
   846 => x"2028676f",
   847 => x"74203078",
   848 => x"2564290a",
   849 => x"00000000",
   850 => x"42797465",
   851 => x"20636865",
   852 => x"636b2066",
   853 => x"61696c65",
   854 => x"64202861",
   855 => x"66746572",
   856 => x"20636163",
   857 => x"68652072",
   858 => x"65667265",
   859 => x"73682920",
   860 => x"61742033",
   861 => x"2028676f",
   862 => x"74203078",
   863 => x"2564290a",
   864 => x"00000000",
   865 => x"43686563",
   866 => x"6b696e67",
   867 => x"206d656d",
   868 => x"6f72792e",
   869 => x"2e2e0a00",
   870 => x"30782564",
   871 => x"20676f6f",
   872 => x"64207265",
   873 => x"6164732c",
   874 => x"20000000",
   875 => x"4572726f",
   876 => x"72206174",
   877 => x"20307825",
   878 => x"642c2065",
   879 => x"78706563",
   880 => x"74656420",
   881 => x"30782564",
   882 => x"2c20676f",
   883 => x"74203078",
   884 => x"25640a00",
   885 => x"42616420",
   886 => x"64617461",
   887 => x"20666f75",
   888 => x"6e642061",
   889 => x"74203078",
   890 => x"25642028",
   891 => x"30782564",
   892 => x"290a0000",
   893 => x"416c6961",
   894 => x"73657320",
   895 => x"666f756e",
   896 => x"64206174",
   897 => x"20307825",
   898 => x"640a0000",
   899 => x"28416c69",
   900 => x"61736573",
   901 => x"2070726f",
   902 => x"6261626c",
   903 => x"79207369",
   904 => x"6d706c79",
   905 => x"20696e64",
   906 => x"69636174",
   907 => x"65207468",
   908 => x"61742052",
   909 => x"414d2069",
   910 => x"7320736d",
   911 => x"616c6c65",
   912 => x"72207468",
   913 => x"616e2036",
   914 => x"34206d65",
   915 => x"67616279",
   916 => x"74657329",
   917 => x"00000000",
   918 => x"53445241",
   919 => x"4d207369",
   920 => x"7a652028",
   921 => x"61737375",
   922 => x"6d696e67",
   923 => x"206e6f20",
   924 => x"61646472",
   925 => x"65737320",
   926 => x"6661756c",
   927 => x"74732920",
   928 => x"69732030",
   929 => x"78256420",
   930 => x"6d656761",
   931 => x"62797465",
   932 => x"730a0000",
   933 => x"46697273",
   934 => x"74207374",
   935 => x"61676520",
   936 => x"73616e69",
   937 => x"74792063",
   938 => x"6865636b",
   939 => x"20706173",
   940 => x"7365642e",
   941 => x"0a000000",
   942 => x"42797465",
   943 => x"20286471",
   944 => x"6d292063",
   945 => x"6865636b",
   946 => x"20706173",
   947 => x"7365640a",
   948 => x"00000000",
   949 => x"41646472",
   950 => x"65737320",
   951 => x"63686563",
   952 => x"6b207061",
   953 => x"73736564",
   954 => x"2e0a0000",
   955 => x"4c465352",
   956 => x"20636865",
   957 => x"636b2070",
   958 => x"61737365",
   959 => x"642e0a00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

