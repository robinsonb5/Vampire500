-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08080f4",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"8a907383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"803d0d91",
    30 => x"3fa0808a",
    31 => x"a0518397",
    32 => x"3f800b80",
    33 => x"0c823d0d",
    34 => x"04fe3d0d",
    35 => x"fea0800b",
    36 => x"86ffe280",
    37 => x"23800b86",
    38 => x"ffe28223",
    39 => x"800b86ff",
    40 => x"e2842380",
    41 => x"0b86ffe2",
    42 => x"8823800b",
    43 => x"86ffe28a",
    44 => x"23907053",
    45 => x"53a0bf51",
    46 => x"80727084",
    47 => x"05540cff",
    48 => x"11517080",
    49 => x"25f238bc",
    50 => x"0b86ffe1",
    51 => x"922381d4",
    52 => x"0b86ffe1",
    53 => x"942380d9",
    54 => x"810b86ff",
    55 => x"e18e23e9",
    56 => x"c10b86ff",
    57 => x"e1902386",
    58 => x"ff0b86ff",
    59 => x"e380239f",
    60 => x"ff0b86ff",
    61 => x"e3822381",
    62 => x"e00b8488",
    63 => x"9023900b",
    64 => x"902c5170",
    65 => x"84889223",
    66 => x"81e20b84",
    67 => x"88942372",
    68 => x"84889623",
    69 => x"ff0b8488",
    70 => x"9823fe0b",
    71 => x"84889a23",
    72 => x"8488900b",
    73 => x"902c5271",
    74 => x"86ffe180",
    75 => x"23848890",
    76 => x"517086ff",
    77 => x"e1822380",
    78 => x"0b86ffe1",
    79 => x"8823fe87",
    80 => x"900b86ff",
    81 => x"e1962380",
    82 => x"0b8488a0",
    83 => x"0c800b84",
    84 => x"88a40c84",
    85 => x"3d0d04f9",
    86 => x"3d0d02a7",
    87 => x"05338488",
    88 => x"a4088488",
    89 => x"a0087184",
    90 => x"b0291190",
    91 => x"1174a029",
    92 => x"19f88011",
    93 => x"08f88412",
    94 => x"08525a5a",
    95 => x"51565a58",
    96 => x"56737334",
    97 => x"73ffb014",
    98 => x"3473fee0",
    99 => x"143473fe",
   100 => x"90143474",
   101 => x"fdc01434",
   102 => x"74fcf014",
   103 => x"3474fca0",
   104 => x"143474fb",
   105 => x"d0143475",
   106 => x"8a2e80de",
   107 => x"38811884",
   108 => x"88a00c84",
   109 => x"88a00880",
   110 => x"d02eb238",
   111 => x"76992e85",
   112 => x"38893d0d",
   113 => x"04900b94",
   114 => x"80115654",
   115 => x"9f9f5374",
   116 => x"70840556",
   117 => x"08747084",
   118 => x"05560cff",
   119 => x"13537280",
   120 => x"25ed3898",
   121 => x"0b8488a4",
   122 => x"0c893d0d",
   123 => x"04811784",
   124 => x"88a40c80",
   125 => x"0b8488a0",
   126 => x"0c8488a4",
   127 => x"08577699",
   128 => x"2e098106",
   129 => x"ffbb38ff",
   130 => x"bc398117",
   131 => x"8488a40c",
   132 => x"8488a408",
   133 => x"57e839f5",
   134 => x"3d0d7d5c",
   135 => x"7b708405",
   136 => x"5d085a80",
   137 => x"5979982a",
   138 => x"7a882b5b",
   139 => x"5877802e",
   140 => x"80f13884",
   141 => x"88a40884",
   142 => x"88a00871",
   143 => x"84b02911",
   144 => x"90117ba0",
   145 => x"2917f880",
   146 => x"1108f884",
   147 => x"1208f888",
   148 => x"13535c5a",
   149 => x"5751565c",
   150 => x"57747434",
   151 => x"74ffb015",
   152 => x"3474fee0",
   153 => x"153474fe",
   154 => x"90153475",
   155 => x"fdc01534",
   156 => x"75fcf015",
   157 => x"3475fca0",
   158 => x"153475fb",
   159 => x"d0153477",
   160 => x"8a2e80f3",
   161 => x"38811b84",
   162 => x"88a00c84",
   163 => x"88a00880",
   164 => x"d02e80c6",
   165 => x"3876992e",
   166 => x"92388119",
   167 => x"59837925",
   168 => x"ff833877",
   169 => x"fef6388d",
   170 => x"3d0d0490",
   171 => x"0b948011",
   172 => x"57559f9f",
   173 => x"54757084",
   174 => x"05570875",
   175 => x"70840557",
   176 => x"0cff1454",
   177 => x"738025ed",
   178 => x"38980b84",
   179 => x"88a40c81",
   180 => x"19598379",
   181 => x"25fece38",
   182 => x"ca398117",
   183 => x"8488a40c",
   184 => x"800b8488",
   185 => x"a00c8488",
   186 => x"a4085776",
   187 => x"992e0981",
   188 => x"06ffa738",
   189 => x"ffb53981",
   190 => x"178488a4",
   191 => x"0c8488a4",
   192 => x"0857e839",
   193 => x"ff3d0d02",
   194 => x"8f053352",
   195 => x"ff840870",
   196 => x"882a7081",
   197 => x"06515151",
   198 => x"70802ef0",
   199 => x"3871ff84",
   200 => x"0c833d0d",
   201 => x"04fe3d0d",
   202 => x"74703352",
   203 => x"5370802e",
   204 => x"a1387052",
   205 => x"811353ff",
   206 => x"84087088",
   207 => x"2a708106",
   208 => x"51515170",
   209 => x"802ef038",
   210 => x"71ff840c",
   211 => x"72335271",
   212 => x"e338843d",
   213 => x"0d04ff3d",
   214 => x"0dff8408",
   215 => x"70892a70",
   216 => x"81065152",
   217 => x"5270802e",
   218 => x"f0387181",
   219 => x"ff06800c",
   220 => x"833d0d04",
   221 => x"ff3d0d02",
   222 => x"8f053352",
   223 => x"ff840870",
   224 => x"882a7081",
   225 => x"06515151",
   226 => x"70802ef0",
   227 => x"3871ff84",
   228 => x"0c833d0d",
   229 => x"04f53d0d",
   230 => x"8e3d7070",
   231 => x"84055208",
   232 => x"a08086f4",
   233 => x"5b555b80",
   234 => x"74708105",
   235 => x"5633755a",
   236 => x"54577277",
   237 => x"2ebe3872",
   238 => x"a52e0981",
   239 => x"0680c538",
   240 => x"77708105",
   241 => x"59335372",
   242 => x"80e42e81",
   243 => x"b6387280",
   244 => x"e42480c6",
   245 => x"387280e3",
   246 => x"2ea13880",
   247 => x"52a55178",
   248 => x"2d805272",
   249 => x"51782d82",
   250 => x"17577770",
   251 => x"81055933",
   252 => x"5372c438",
   253 => x"76800c8d",
   254 => x"3d0d047a",
   255 => x"841c8312",
   256 => x"33555c56",
   257 => x"80527251",
   258 => x"782d8117",
   259 => x"78708105",
   260 => x"5a335457",
   261 => x"72ffa038",
   262 => x"db397280",
   263 => x"f32e0981",
   264 => x"06ffb838",
   265 => x"7a841c71",
   266 => x"08585c54",
   267 => x"8076335b",
   268 => x"5579752e",
   269 => x"8d388115",
   270 => x"70177033",
   271 => x"555b5572",
   272 => x"f538ff15",
   273 => x"54807525",
   274 => x"ffa03875",
   275 => x"70810557",
   276 => x"33538052",
   277 => x"7251782d",
   278 => x"811774ff",
   279 => x"16565657",
   280 => x"807525ff",
   281 => x"85387570",
   282 => x"81055733",
   283 => x"53805272",
   284 => x"51782d81",
   285 => x"1774ff16",
   286 => x"56565774",
   287 => x"8024cc38",
   288 => x"fee8397a",
   289 => x"841c7108",
   290 => x"8488f80b",
   291 => x"8488a854",
   292 => x"5d565c55",
   293 => x"80567376",
   294 => x"2e098106",
   295 => x"b838b00b",
   296 => x"8488a834",
   297 => x"811555ff",
   298 => x"15557433",
   299 => x"7a708105",
   300 => x"5c348116",
   301 => x"56748488",
   302 => x"a82e0981",
   303 => x"06e93880",
   304 => x"7a347584",
   305 => x"88f80bff",
   306 => x"12565755",
   307 => x"748024fe",
   308 => x"fa38fe96",
   309 => x"39738f06",
   310 => x"a08098b0",
   311 => x"05537233",
   312 => x"75708105",
   313 => x"57347384",
   314 => x"2a5473e9",
   315 => x"38748488",
   316 => x"a82ecc38",
   317 => x"ff155574",
   318 => x"337a7081",
   319 => x"055c3481",
   320 => x"16567484",
   321 => x"88a82eff",
   322 => x"b638ff9b",
   323 => x"39000000",
   324 => x"00ffffff",
   325 => x"ff00ffff",
   326 => x"ffff00ff",
   327 => x"ffffff00",
   328 => x"48656c6c",
   329 => x"6f2c2077",
   330 => x"6f726c64",
   331 => x"210a0000",
   332 => x"00000000",
   333 => x"00000000",
   334 => x"18181818",
   335 => x"18001800",
   336 => x"6c6c0000",
   337 => x"00000000",
   338 => x"6c6cfe6c",
   339 => x"fe6c6c00",
   340 => x"183e603c",
   341 => x"067c1800",
   342 => x"0066acd8",
   343 => x"366acc00",
   344 => x"386c6876",
   345 => x"dcce7b00",
   346 => x"18183000",
   347 => x"00000000",
   348 => x"0c183030",
   349 => x"30180c00",
   350 => x"30180c0c",
   351 => x"0c183000",
   352 => x"00663cff",
   353 => x"3c660000",
   354 => x"0018187e",
   355 => x"18180000",
   356 => x"00000000",
   357 => x"00181830",
   358 => x"0000007e",
   359 => x"00000000",
   360 => x"00000000",
   361 => x"00181800",
   362 => x"03060c18",
   363 => x"3060c000",
   364 => x"3c666e7e",
   365 => x"76663c00",
   366 => x"18387818",
   367 => x"18181800",
   368 => x"3c66060c",
   369 => x"18307e00",
   370 => x"3c66061c",
   371 => x"06663c00",
   372 => x"1c3c6ccc",
   373 => x"fe0c0c00",
   374 => x"7e607c06",
   375 => x"06663c00",
   376 => x"1c30607c",
   377 => x"66663c00",
   378 => x"7e06060c",
   379 => x"18181800",
   380 => x"3c66663c",
   381 => x"66663c00",
   382 => x"3c66663e",
   383 => x"060c3800",
   384 => x"00181800",
   385 => x"00181800",
   386 => x"00181800",
   387 => x"00181830",
   388 => x"00061860",
   389 => x"18060000",
   390 => x"00007e00",
   391 => x"7e000000",
   392 => x"00601806",
   393 => x"18600000",
   394 => x"3c66060c",
   395 => x"18001800",
   396 => x"7cc6ded6",
   397 => x"dec07800",
   398 => x"3c66667e",
   399 => x"66666600",
   400 => x"7c66667c",
   401 => x"66667c00",
   402 => x"1e306060",
   403 => x"60301e00",
   404 => x"786c6666",
   405 => x"666c7800",
   406 => x"7e606078",
   407 => x"60607e00",
   408 => x"7e606078",
   409 => x"60606000",
   410 => x"3c66606e",
   411 => x"66663e00",
   412 => x"6666667e",
   413 => x"66666600",
   414 => x"3c181818",
   415 => x"18183c00",
   416 => x"06060606",
   417 => x"06663c00",
   418 => x"c6ccd8f0",
   419 => x"d8ccc600",
   420 => x"60606060",
   421 => x"60607e00",
   422 => x"c6eefed6",
   423 => x"c6c6c600",
   424 => x"c6e6f6de",
   425 => x"cec6c600",
   426 => x"3c666666",
   427 => x"66663c00",
   428 => x"7c66667c",
   429 => x"60606000",
   430 => x"78cccccc",
   431 => x"ccdc7e00",
   432 => x"7c66667c",
   433 => x"6c666600",
   434 => x"3c66703c",
   435 => x"0e663c00",
   436 => x"7e181818",
   437 => x"18181800",
   438 => x"66666666",
   439 => x"66663c00",
   440 => x"66666666",
   441 => x"3c3c1800",
   442 => x"c6c6c6d6",
   443 => x"feeec600",
   444 => x"c3663c18",
   445 => x"3c66c300",
   446 => x"c3663c18",
   447 => x"18181800",
   448 => x"fe0c1830",
   449 => x"60c0fe00",
   450 => x"3c303030",
   451 => x"30303c00",
   452 => x"c0603018",
   453 => x"0c060300",
   454 => x"3c0c0c0c",
   455 => x"0c0c3c00",
   456 => x"10386cc6",
   457 => x"00000000",
   458 => x"00000000",
   459 => x"000000fe",
   460 => x"18180c00",
   461 => x"00000000",
   462 => x"00003c06",
   463 => x"3e663e00",
   464 => x"60607c66",
   465 => x"66667c00",
   466 => x"00003c60",
   467 => x"60603c00",
   468 => x"06063e66",
   469 => x"66663e00",
   470 => x"00003c66",
   471 => x"7e603c00",
   472 => x"1c307c30",
   473 => x"30303000",
   474 => x"00003e66",
   475 => x"663e063c",
   476 => x"60607c66",
   477 => x"66666600",
   478 => x"18001818",
   479 => x"18180c00",
   480 => x"0c000c0c",
   481 => x"0c0c0c78",
   482 => x"6060666c",
   483 => x"786c6600",
   484 => x"18181818",
   485 => x"18180c00",
   486 => x"0000ecfe",
   487 => x"d6c6c600",
   488 => x"00007c66",
   489 => x"66666600",
   490 => x"00003c66",
   491 => x"66663c00",
   492 => x"00007c66",
   493 => x"667c6060",
   494 => x"00003e66",
   495 => x"663e0606",
   496 => x"00007c66",
   497 => x"60606000",
   498 => x"00003c60",
   499 => x"3c067c00",
   500 => x"30307c30",
   501 => x"30301c00",
   502 => x"00006666",
   503 => x"66663e00",
   504 => x"00006666",
   505 => x"663c1800",
   506 => x"0000c6c6",
   507 => x"d6fe6c00",
   508 => x"0000c66c",
   509 => x"386cc600",
   510 => x"00006666",
   511 => x"663c1830",
   512 => x"00007e0c",
   513 => x"18307e00",
   514 => x"0e181870",
   515 => x"18180e00",
   516 => x"18181818",
   517 => x"18181800",
   518 => x"7018180e",
   519 => x"18187000",
   520 => x"729c0000",
   521 => x"00000000",
   522 => x"fefefefe",
   523 => x"fefefe00",
   524 => x"00000000",
   525 => x"00000000",
   526 => x"00000000",
   527 => x"00000000",
   528 => x"00000000",
   529 => x"00000000",
   530 => x"00000000",
   531 => x"00000000",
   532 => x"00000000",
   533 => x"00000000",
   534 => x"00000000",
   535 => x"00000000",
   536 => x"00000000",
   537 => x"00000000",
   538 => x"00000000",
   539 => x"00000000",
   540 => x"00000000",
   541 => x"00000000",
   542 => x"00000000",
   543 => x"00000000",
   544 => x"00000000",
   545 => x"00000000",
   546 => x"00000000",
   547 => x"00000000",
   548 => x"00000000",
   549 => x"00000000",
   550 => x"00000000",
   551 => x"00000000",
   552 => x"00000000",
   553 => x"00000000",
   554 => x"00000000",
   555 => x"00000000",
   556 => x"00000000",
   557 => x"00000000",
   558 => x"00000000",
   559 => x"00000000",
   560 => x"00000000",
   561 => x"00000000",
   562 => x"00000000",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"30313233",
   781 => x"34353637",
   782 => x"38394142",
   783 => x"43444546",
   784 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

