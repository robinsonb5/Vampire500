-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VampireDiag_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VampireDiag_ROM;

architecture arch of VampireDiag_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"a08081a3",
     1 => x"04000000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"89e87383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040000",
    29 => x"02ec050d",
    30 => x"76548755",
    31 => x"739c2a74",
    32 => x"842bb712",
    33 => x"55555271",
    34 => x"89248438",
    35 => x"b0125372",
    36 => x"51a08085",
    37 => x"ea2dff15",
    38 => x"55748025",
    39 => x"df380294",
    40 => x"050d0402",
    41 => x"e4050d83",
    42 => x"0b85ffc4",
    43 => x"8134fc0b",
    44 => x"85ffc081",
    45 => x"34a08083",
    46 => x"a62d87f0",
    47 => x"80802287",
    48 => x"f0808022",
    49 => x"70902b70",
    50 => x"902c8422",
    51 => x"52525254",
    52 => x"52800b9e",
    53 => x"800a2270",
    54 => x"902b7090",
    55 => x"2c595656",
    56 => x"5772762e",
    57 => x"09810699",
    58 => x"38811784",
    59 => x"229e800a",
    60 => x"2270902b",
    61 => x"70902c5a",
    62 => x"57575357",
    63 => x"72762ee9",
    64 => x"3887f080",
    65 => x"8422a080",
    66 => x"89f85252",
    67 => x"a08087d1",
    68 => x"2d725487",
    69 => x"55739c2a",
    70 => x"74842bb7",
    71 => x"12555552",
    72 => x"71892484",
    73 => x"38b01253",
    74 => x"7251a080",
    75 => x"85ea2dff",
    76 => x"15557480",
    77 => x"25df38a0",
    78 => x"808a8451",
    79 => x"a08087d1",
    80 => x"2d765487",
    81 => x"55739c2a",
    82 => x"74842bb7",
    83 => x"12555552",
    84 => x"71892484",
    85 => x"38b01253",
    86 => x"7251a080",
    87 => x"85ea2dff",
    88 => x"15557480",
    89 => x"25df38a0",
    90 => x"808a9451",
    91 => x"a08087d1",
    92 => x"2da0808a",
    93 => x"a851a080",
    94 => x"87d12d75",
    95 => x"54875573",
    96 => x"9c2a7484",
    97 => x"2bb71255",
    98 => x"55527189",
    99 => x"248438b0",
   100 => x"12537251",
   101 => x"a08085ea",
   102 => x"2dff1555",
   103 => x"748025df",
   104 => x"38a08083",
   105 => x"a10402f4",
   106 => x"050dfea0",
   107 => x"800b86ff",
   108 => x"e2802380",
   109 => x"0b86ffe2",
   110 => x"8223800b",
   111 => x"86ffe284",
   112 => x"23800b86",
   113 => x"ffe28823",
   114 => x"800b86ff",
   115 => x"e28a2390",
   116 => x"705353a0",
   117 => x"bf518072",
   118 => x"70840554",
   119 => x"0cff1151",
   120 => x"708025f2",
   121 => x"38bc0b86",
   122 => x"ffe19223",
   123 => x"81d40b86",
   124 => x"ffe19423",
   125 => x"80d9810b",
   126 => x"86ffe18e",
   127 => x"23e9c10b",
   128 => x"86ffe190",
   129 => x"2386ff0b",
   130 => x"86ffe380",
   131 => x"239fff0b",
   132 => x"86ffe382",
   133 => x"2381e00b",
   134 => x"84889023",
   135 => x"900b902c",
   136 => x"51708488",
   137 => x"922381e2",
   138 => x"0b848894",
   139 => x"23728488",
   140 => x"9623ff0b",
   141 => x"84889823",
   142 => x"fe0b8488",
   143 => x"9a238488",
   144 => x"900b902c",
   145 => x"527186ff",
   146 => x"e1802384",
   147 => x"88905170",
   148 => x"86ffe182",
   149 => x"23800b86",
   150 => x"ffe18823",
   151 => x"fe87900b",
   152 => x"86ffe196",
   153 => x"23800b84",
   154 => x"88a00c80",
   155 => x"0b8488a4",
   156 => x"0c028c05",
   157 => x"0d0402f8",
   158 => x"050d8488",
   159 => x"a4081010",
   160 => x"8488a408",
   161 => x"05709029",
   162 => x"8488a008",
   163 => x"0584c011",
   164 => x"51525280",
   165 => x"52717134",
   166 => x"71811234",
   167 => x"71821234",
   168 => x"71831234",
   169 => x"80d01181",
   170 => x"13535181",
   171 => x"ff7225e5",
   172 => x"38028805",
   173 => x"0d0402f4",
   174 => x"050d9053",
   175 => x"a0bf5272",
   176 => x"84147108",
   177 => x"8105720c",
   178 => x"ff145454",
   179 => x"51807224",
   180 => x"e9387284",
   181 => x"14710881",
   182 => x"05720cff",
   183 => x"14545451",
   184 => x"718025db",
   185 => x"38a08085",
   186 => x"ba0402e8",
   187 => x"050d7756",
   188 => x"9f762581",
   189 => x"8d388488",
   190 => x"a4087010",
   191 => x"10117081",
   192 => x"80298488",
   193 => x"a0080584",
   194 => x"c0117910",
   195 => x"1010a080",
   196 => x"88c00570",
   197 => x"70840552",
   198 => x"08710852",
   199 => x"54555154",
   200 => x"55557072",
   201 => x"3470882c",
   202 => x"5372ffb0",
   203 => x"13347090",
   204 => x"2c5372fe",
   205 => x"e0133470",
   206 => x"982c5170",
   207 => x"fe901334",
   208 => x"73fdc013",
   209 => x"3473882c",
   210 => x"5372fcf0",
   211 => x"13347390",
   212 => x"2c5170fc",
   213 => x"a0133473",
   214 => x"982c5473",
   215 => x"fbd01334",
   216 => x"758a2eab",
   217 => x"388488a0",
   218 => x"08810584",
   219 => x"88a00c84",
   220 => x"88a00880",
   221 => x"d02e9838",
   222 => x"74992eac",
   223 => x"38029805",
   224 => x"0d048488",
   225 => x"a4085575",
   226 => x"8a2e0981",
   227 => x"06d73881",
   228 => x"158488a4",
   229 => x"0c800b84",
   230 => x"88a00c84",
   231 => x"88a40855",
   232 => x"74992e09",
   233 => x"8106d638",
   234 => x"900b9480",
   235 => x"1154529f",
   236 => x"9f517270",
   237 => x"84055408",
   238 => x"72708405",
   239 => x"540cff11",
   240 => x"51708025",
   241 => x"ed38980b",
   242 => x"8488a40c",
   243 => x"0298050d",
   244 => x"0402dc05",
   245 => x"0d7a5877",
   246 => x"70840559",
   247 => x"08578059",
   248 => x"76982a77",
   249 => x"882b5856",
   250 => x"75802e81",
   251 => x"9b389f76",
   252 => x"25819a38",
   253 => x"8488a408",
   254 => x"70101011",
   255 => x"70818029",
   256 => x"8488a008",
   257 => x"0584c011",
   258 => x"79101010",
   259 => x"a08088c0",
   260 => x"05707084",
   261 => x"05520871",
   262 => x"08525455",
   263 => x"51545555",
   264 => x"70723470",
   265 => x"882c5372",
   266 => x"ffb01334",
   267 => x"70902c53",
   268 => x"72fee013",
   269 => x"3470982c",
   270 => x"5170fe90",
   271 => x"133473fd",
   272 => x"c0133473",
   273 => x"882c5372",
   274 => x"fcf01334",
   275 => x"73902c51",
   276 => x"70fca013",
   277 => x"3473982c",
   278 => x"5473fbd0",
   279 => x"1334758a",
   280 => x"2eb83884",
   281 => x"88a00881",
   282 => x"058488a0",
   283 => x"0c8488a0",
   284 => x"0880d02e",
   285 => x"a5387499",
   286 => x"2eb93881",
   287 => x"19598379",
   288 => x"25fedd38",
   289 => x"75fed038",
   290 => x"02a4050d",
   291 => x"048488a4",
   292 => x"0855758a",
   293 => x"2e098106",
   294 => x"ca388115",
   295 => x"8488a40c",
   296 => x"800b8488",
   297 => x"a00c8488",
   298 => x"a4085574",
   299 => x"992e0981",
   300 => x"06c93890",
   301 => x"0b948011",
   302 => x"54529f9f",
   303 => x"51727084",
   304 => x"05540872",
   305 => x"70840554",
   306 => x"0cff1151",
   307 => x"708025ed",
   308 => x"38980b84",
   309 => x"88a40c81",
   310 => x"19598379",
   311 => x"25fe8138",
   312 => x"a0808984",
   313 => x"04000000",
   314 => x"00ffffff",
   315 => x"ff00ffff",
   316 => x"ffff00ff",
   317 => x"ffffff00",
   318 => x"53686164",
   319 => x"6f77206f",
   320 => x"66200000",
   321 => x"20706572",
   322 => x"73697374",
   323 => x"65642066",
   324 => x"6f722000",
   325 => x"20636f6e",
   326 => x"73656375",
   327 => x"74697665",
   328 => x"20726561",
   329 => x"64730a00",
   330 => x"456e6469",
   331 => x"6e672077",
   332 => x"69746820",
   333 => x"61207265",
   334 => x"6164206f",
   335 => x"66200000",
   336 => x"00000000",
   337 => x"00000000",
   338 => x"18181818",
   339 => x"18001800",
   340 => x"6c6c0000",
   341 => x"00000000",
   342 => x"6c6cfe6c",
   343 => x"fe6c6c00",
   344 => x"183e603c",
   345 => x"067c1800",
   346 => x"0066acd8",
   347 => x"366acc00",
   348 => x"386c6876",
   349 => x"dcce7b00",
   350 => x"18183000",
   351 => x"00000000",
   352 => x"0c183030",
   353 => x"30180c00",
   354 => x"30180c0c",
   355 => x"0c183000",
   356 => x"00663cff",
   357 => x"3c660000",
   358 => x"0018187e",
   359 => x"18180000",
   360 => x"00000000",
   361 => x"00181830",
   362 => x"0000007e",
   363 => x"00000000",
   364 => x"00000000",
   365 => x"00181800",
   366 => x"03060c18",
   367 => x"3060c000",
   368 => x"3c666e7e",
   369 => x"76663c00",
   370 => x"18387818",
   371 => x"18181800",
   372 => x"3c66060c",
   373 => x"18307e00",
   374 => x"3c66061c",
   375 => x"06663c00",
   376 => x"1c3c6ccc",
   377 => x"fe0c0c00",
   378 => x"7e607c06",
   379 => x"06663c00",
   380 => x"1c30607c",
   381 => x"66663c00",
   382 => x"7e06060c",
   383 => x"18181800",
   384 => x"3c66663c",
   385 => x"66663c00",
   386 => x"3c66663e",
   387 => x"060c3800",
   388 => x"00181800",
   389 => x"00181800",
   390 => x"00181800",
   391 => x"00181830",
   392 => x"00061860",
   393 => x"18060000",
   394 => x"00007e00",
   395 => x"7e000000",
   396 => x"00601806",
   397 => x"18600000",
   398 => x"3c66060c",
   399 => x"18001800",
   400 => x"7cc6ded6",
   401 => x"dec07800",
   402 => x"3c66667e",
   403 => x"66666600",
   404 => x"7c66667c",
   405 => x"66667c00",
   406 => x"1e306060",
   407 => x"60301e00",
   408 => x"786c6666",
   409 => x"666c7800",
   410 => x"7e606078",
   411 => x"60607e00",
   412 => x"7e606078",
   413 => x"60606000",
   414 => x"3c66606e",
   415 => x"66663e00",
   416 => x"6666667e",
   417 => x"66666600",
   418 => x"3c181818",
   419 => x"18183c00",
   420 => x"06060606",
   421 => x"06663c00",
   422 => x"c6ccd8f0",
   423 => x"d8ccc600",
   424 => x"60606060",
   425 => x"60607e00",
   426 => x"c6eefed6",
   427 => x"c6c6c600",
   428 => x"c6e6f6de",
   429 => x"cec6c600",
   430 => x"3c666666",
   431 => x"66663c00",
   432 => x"7c66667c",
   433 => x"60606000",
   434 => x"78cccccc",
   435 => x"ccdc7e00",
   436 => x"7c66667c",
   437 => x"6c666600",
   438 => x"3c66703c",
   439 => x"0e663c00",
   440 => x"7e181818",
   441 => x"18181800",
   442 => x"66666666",
   443 => x"66663c00",
   444 => x"66666666",
   445 => x"3c3c1800",
   446 => x"c6c6c6d6",
   447 => x"feeec600",
   448 => x"c3663c18",
   449 => x"3c66c300",
   450 => x"c3663c18",
   451 => x"18181800",
   452 => x"fe0c1830",
   453 => x"60c0fe00",
   454 => x"3c303030",
   455 => x"30303c00",
   456 => x"c0603018",
   457 => x"0c060300",
   458 => x"3c0c0c0c",
   459 => x"0c0c3c00",
   460 => x"10386cc6",
   461 => x"00000000",
   462 => x"00000000",
   463 => x"000000fe",
   464 => x"18180c00",
   465 => x"00000000",
   466 => x"00003c06",
   467 => x"3e663e00",
   468 => x"60607c66",
   469 => x"66667c00",
   470 => x"00003c60",
   471 => x"60603c00",
   472 => x"06063e66",
   473 => x"66663e00",
   474 => x"00003c66",
   475 => x"7e603c00",
   476 => x"1c307c30",
   477 => x"30303000",
   478 => x"00003e66",
   479 => x"663e063c",
   480 => x"60607c66",
   481 => x"66666600",
   482 => x"18001818",
   483 => x"18180c00",
   484 => x"0c000c0c",
   485 => x"0c0c0c78",
   486 => x"6060666c",
   487 => x"786c6600",
   488 => x"18181818",
   489 => x"18180c00",
   490 => x"0000ecfe",
   491 => x"d6c6c600",
   492 => x"00007c66",
   493 => x"66666600",
   494 => x"00003c66",
   495 => x"66663c00",
   496 => x"00007c66",
   497 => x"667c6060",
   498 => x"00003e66",
   499 => x"663e0606",
   500 => x"00007c66",
   501 => x"60606000",
   502 => x"00003c60",
   503 => x"3c067c00",
   504 => x"30307c30",
   505 => x"30301c00",
   506 => x"00006666",
   507 => x"66663e00",
   508 => x"00006666",
   509 => x"663c1800",
   510 => x"0000c6c6",
   511 => x"d6fe6c00",
   512 => x"0000c66c",
   513 => x"386cc600",
   514 => x"00006666",
   515 => x"663c1830",
   516 => x"00007e0c",
   517 => x"18307e00",
   518 => x"0e181870",
   519 => x"18180e00",
   520 => x"18181818",
   521 => x"18181800",
   522 => x"7018180e",
   523 => x"18187000",
   524 => x"729c0000",
   525 => x"00000000",
   526 => x"fefefefe",
   527 => x"fefefe00",
   528 => x"00000000",
   529 => x"00000000",
   530 => x"00000000",
   531 => x"00000000",
   532 => x"00000000",
   533 => x"00000000",
   534 => x"00000000",
   535 => x"00000000",
   536 => x"00000000",
   537 => x"00000000",
   538 => x"00000000",
   539 => x"00000000",
   540 => x"00000000",
   541 => x"00000000",
   542 => x"00000000",
   543 => x"00000000",
   544 => x"00000000",
   545 => x"00000000",
   546 => x"00000000",
   547 => x"00000000",
   548 => x"00000000",
   549 => x"00000000",
   550 => x"00000000",
   551 => x"00000000",
   552 => x"00000000",
   553 => x"00000000",
   554 => x"00000000",
   555 => x"00000000",
   556 => x"00000000",
   557 => x"00000000",
   558 => x"00000000",
   559 => x"00000000",
   560 => x"00000000",
   561 => x"00000000",
   562 => x"00000000",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000000",
   592 => x"00000000",
   593 => x"00000000",
   594 => x"00000000",
   595 => x"00000000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

