-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"f2040000",
     2 => x"800b810b",
     3 => x"ff8c0c04",
     4 => x"0b0b0ba0",
     5 => x"80809d0b",
     6 => x"810bff8c",
     7 => x"0c700471",
     8 => x"fd060872",
     9 => x"83060981",
    10 => x"05820583",
    11 => x"2b2a83ff",
    12 => x"ff065204",
    13 => x"71fc0608",
    14 => x"72830609",
    15 => x"81058305",
    16 => x"1010102a",
    17 => x"81ff0652",
    18 => x"0471fc06",
    19 => x"080ba080",
    20 => x"93c47383",
    21 => x"06101005",
    22 => x"08067381",
    23 => x"ff067383",
    24 => x"06098105",
    25 => x"83051010",
    26 => x"102b0772",
    27 => x"fc060c51",
    28 => x"51040ba0",
    29 => x"8080fd0b",
    30 => x"a08092da",
    31 => x"040ba080",
    32 => x"80fd0402",
    33 => x"f8050d02",
    34 => x"8f05a080",
    35 => x"80b42d52",
    36 => x"ff840870",
    37 => x"882a7081",
    38 => x"06515151",
    39 => x"70802ef0",
    40 => x"3871ff84",
    41 => x"0c028805",
    42 => x"0d0402f4",
    43 => x"050d7453",
    44 => x"72a08080",
    45 => x"b42d7081",
    46 => x"ff065252",
    47 => x"70802ea3",
    48 => x"387181ff",
    49 => x"06811454",
    50 => x"52ff8408",
    51 => x"70882a70",
    52 => x"81065151",
    53 => x"5170802e",
    54 => x"f03871ff",
    55 => x"840ca080",
    56 => x"81b00402",
    57 => x"8c050d04",
    58 => x"02f8050d",
    59 => x"028f05a0",
    60 => x"8080b42d",
    61 => x"52ff8408",
    62 => x"70882a70",
    63 => x"81065151",
    64 => x"5170802e",
    65 => x"f03871ff",
    66 => x"840c0288",
    67 => x"050d0402",
    68 => x"d0050d02",
    69 => x"b405a080",
    70 => x"81e87170",
    71 => x"84055308",
    72 => x"5c5c5880",
    73 => x"7a708105",
    74 => x"5ca08080",
    75 => x"b42d5459",
    76 => x"72792e82",
    77 => x"cc3872a5",
    78 => x"2e098106",
    79 => x"82ab3879",
    80 => x"7081055b",
    81 => x"a08080b4",
    82 => x"2d537280",
    83 => x"e42e9f38",
    84 => x"7280e424",
    85 => x"8d387280",
    86 => x"e32e81c4",
    87 => x"38a08084",
    88 => x"b2047280",
    89 => x"f32e818d",
    90 => x"38a08084",
    91 => x"b2047784",
    92 => x"19710883",
    93 => x"ffe0e00b",
    94 => x"83ffe090",
    95 => x"595a5659",
    96 => x"53805673",
    97 => x"762e0981",
    98 => x"069538b0",
    99 => x"0b83ffe0",
   100 => x"900ba080",
   101 => x"80c92d81",
   102 => x"1555a080",
   103 => x"83c70473",
   104 => x"8f06a080",
   105 => x"93d40553",
   106 => x"72a08080",
   107 => x"b42d7570",
   108 => x"810557a0",
   109 => x"8080c92d",
   110 => x"73842a54",
   111 => x"73e13874",
   112 => x"83ffe090",
   113 => x"2e9c38ff",
   114 => x"155574a0",
   115 => x"8080b42d",
   116 => x"77708105",
   117 => x"59a08080",
   118 => x"c92d8116",
   119 => x"56a08083",
   120 => x"bf048077",
   121 => x"a08080c9",
   122 => x"2d7583ff",
   123 => x"e0e05654",
   124 => x"a08084c6",
   125 => x"04778419",
   126 => x"71085759",
   127 => x"538075a0",
   128 => x"8080b42d",
   129 => x"54547274",
   130 => x"2ebc3881",
   131 => x"14701670",
   132 => x"a08080b4",
   133 => x"2d515454",
   134 => x"72f138a0",
   135 => x"8084c604",
   136 => x"77841983",
   137 => x"12a08080",
   138 => x"b42d5259",
   139 => x"53a08084",
   140 => x"e9048052",
   141 => x"a5517a2d",
   142 => x"80527251",
   143 => x"7a2d8219",
   144 => x"59a08084",
   145 => x"f20473ff",
   146 => x"15555380",
   147 => x"7325a338",
   148 => x"74708105",
   149 => x"56a08080",
   150 => x"b42d5380",
   151 => x"5272517a",
   152 => x"2d811959",
   153 => x"a08084c6",
   154 => x"04805272",
   155 => x"517a2d81",
   156 => x"19597970",
   157 => x"81055ba0",
   158 => x"8080b42d",
   159 => x"5372fdb6",
   160 => x"387883ff",
   161 => x"e0800c02",
   162 => x"b0050d04",
   163 => x"02f4050d",
   164 => x"74767181",
   165 => x"ff06c80c",
   166 => x"535383ff",
   167 => x"e1a00885",
   168 => x"3871892b",
   169 => x"5271982a",
   170 => x"c80c7190",
   171 => x"2a7081ff",
   172 => x"06c80c51",
   173 => x"71882a70",
   174 => x"81ff06c8",
   175 => x"0c517181",
   176 => x"ff06c80c",
   177 => x"72902a70",
   178 => x"81ff06c8",
   179 => x"0c51c808",
   180 => x"7081ff06",
   181 => x"515182b8",
   182 => x"bf527081",
   183 => x"ff2e0981",
   184 => x"06943881",
   185 => x"ff0bc80c",
   186 => x"c8087081",
   187 => x"ff06ff14",
   188 => x"54515171",
   189 => x"e5387083",
   190 => x"ffe0800c",
   191 => x"028c050d",
   192 => x"0402fc05",
   193 => x"0d81c751",
   194 => x"81ff0bc8",
   195 => x"0cff1151",
   196 => x"708025f4",
   197 => x"38028405",
   198 => x"0d0402f0",
   199 => x"050da080",
   200 => x"86812d81",
   201 => x"9c9f5380",
   202 => x"5287fc80",
   203 => x"f751a080",
   204 => x"858c2d83",
   205 => x"ffe08008",
   206 => x"5483ffe0",
   207 => x"8008812e",
   208 => x"098106ab",
   209 => x"3881ff0b",
   210 => x"c80c820a",
   211 => x"52849c80",
   212 => x"e951a080",
   213 => x"858c2d83",
   214 => x"ffe08008",
   215 => x"8d3881ff",
   216 => x"0bc80c73",
   217 => x"53a08086",
   218 => x"f604a080",
   219 => x"86812dff",
   220 => x"135372ff",
   221 => x"b2387283",
   222 => x"ffe0800c",
   223 => x"0290050d",
   224 => x"0402f405",
   225 => x"0d81ff0b",
   226 => x"c80c9353",
   227 => x"805287fc",
   228 => x"80c151a0",
   229 => x"80858c2d",
   230 => x"83ffe080",
   231 => x"088d3881",
   232 => x"ff0bc80c",
   233 => x"8153a080",
   234 => x"87b604a0",
   235 => x"8086812d",
   236 => x"ff135372",
   237 => x"d7387283",
   238 => x"ffe0800c",
   239 => x"028c050d",
   240 => x"0402f005",
   241 => x"0da08086",
   242 => x"812d83aa",
   243 => x"52849c80",
   244 => x"c851a080",
   245 => x"858c2d83",
   246 => x"ffe08008",
   247 => x"812e0981",
   248 => x"068e38cc",
   249 => x"0883ffff",
   250 => x"06537283",
   251 => x"aa2ea338",
   252 => x"a0808781",
   253 => x"2da08088",
   254 => x"8b048154",
   255 => x"a08089a2",
   256 => x"04a08093",
   257 => x"e851a080",
   258 => x"828f2d80",
   259 => x"54a08089",
   260 => x"a20481ff",
   261 => x"0bc80cb1",
   262 => x"53a08086",
   263 => x"9a2d83ff",
   264 => x"e0800880",
   265 => x"2e80e238",
   266 => x"805287fc",
   267 => x"80fa51a0",
   268 => x"80858c2d",
   269 => x"83ffe080",
   270 => x"08bf3883",
   271 => x"ffe08008",
   272 => x"52a08094",
   273 => x"8451a080",
   274 => x"828f2d81",
   275 => x"ff0bc80c",
   276 => x"c80881ff",
   277 => x"067053a0",
   278 => x"80949052",
   279 => x"54a08082",
   280 => x"8f2dcc08",
   281 => x"74862a70",
   282 => x"81067057",
   283 => x"51515372",
   284 => x"802eaf38",
   285 => x"a08087fa",
   286 => x"0483ffe0",
   287 => x"800852a0",
   288 => x"80948451",
   289 => x"a080828f",
   290 => x"2d72822e",
   291 => x"fef338ff",
   292 => x"135372ff",
   293 => x"8438a080",
   294 => x"94a051a0",
   295 => x"8081aa2d",
   296 => x"72547383",
   297 => x"ffe0800c",
   298 => x"0290050d",
   299 => x"0402f405",
   300 => x"0d810b83",
   301 => x"ffe1a00c",
   302 => x"c408708f",
   303 => x"2a708106",
   304 => x"51515372",
   305 => x"f33872c4",
   306 => x"0ca08086",
   307 => x"812dc408",
   308 => x"708f2a70",
   309 => x"81065151",
   310 => x"5372f338",
   311 => x"810bc40c",
   312 => x"87538052",
   313 => x"84d480c0",
   314 => x"51a08085",
   315 => x"8c2d83ff",
   316 => x"e0800881",
   317 => x"2e098106",
   318 => x"873883ff",
   319 => x"e0800853",
   320 => x"a08094b8",
   321 => x"51a08081",
   322 => x"aa2d7282",
   323 => x"2e098106",
   324 => x"9238a080",
   325 => x"94cc51a0",
   326 => x"8081aa2d",
   327 => x"8053a080",
   328 => x"8b9304ff",
   329 => x"135372ff",
   330 => x"b938a080",
   331 => x"94ec51a0",
   332 => x"8081aa2d",
   333 => x"a08087c1",
   334 => x"2d83ffe0",
   335 => x"800883ff",
   336 => x"e1a00c83",
   337 => x"ffe08008",
   338 => x"802e8b38",
   339 => x"a0809588",
   340 => x"51a08081",
   341 => x"aa2da080",
   342 => x"959c51a0",
   343 => x"8081aa2d",
   344 => x"815287fc",
   345 => x"80d051a0",
   346 => x"80858c2d",
   347 => x"81ff0bc8",
   348 => x"0cc40870",
   349 => x"8f2a7081",
   350 => x"06515153",
   351 => x"72f33872",
   352 => x"c40c81ff",
   353 => x"0bc80ca0",
   354 => x"8095ac51",
   355 => x"a08081aa",
   356 => x"2d815372",
   357 => x"83ffe080",
   358 => x"0c028c05",
   359 => x"0d04800b",
   360 => x"83ffe080",
   361 => x"0c0402e0",
   362 => x"050d797b",
   363 => x"57578058",
   364 => x"c408708f",
   365 => x"2a708106",
   366 => x"51515473",
   367 => x"f3388281",
   368 => x"0bc40c81",
   369 => x"ff0bc80c",
   370 => x"765287fc",
   371 => x"80d151a0",
   372 => x"80858c2d",
   373 => x"80dbc6df",
   374 => x"5583ffe0",
   375 => x"8008802e",
   376 => x"983883ff",
   377 => x"e0800853",
   378 => x"7652a080",
   379 => x"95b851a0",
   380 => x"80828f2d",
   381 => x"a0808cc5",
   382 => x"0481ff0b",
   383 => x"c80cc808",
   384 => x"7081ff06",
   385 => x"51547381",
   386 => x"fe2e0981",
   387 => x"069b3880",
   388 => x"ff55cc08",
   389 => x"76708405",
   390 => x"580cff15",
   391 => x"55748025",
   392 => x"f1388158",
   393 => x"a0808caf",
   394 => x"04ff1555",
   395 => x"74cb3881",
   396 => x"ff0bc80c",
   397 => x"c408708f",
   398 => x"2a708106",
   399 => x"51515473",
   400 => x"f33873c4",
   401 => x"0c7783ff",
   402 => x"e0800c02",
   403 => x"a0050d04",
   404 => x"02f4050d",
   405 => x"7470882a",
   406 => x"83fe8006",
   407 => x"7072982a",
   408 => x"0772882b",
   409 => x"87fc8080",
   410 => x"0673982b",
   411 => x"81f00a06",
   412 => x"71730707",
   413 => x"83ffe080",
   414 => x"0c565153",
   415 => x"51028c05",
   416 => x"0d0402f4",
   417 => x"050d0292",
   418 => x"05227088",
   419 => x"2a71882b",
   420 => x"077083ff",
   421 => x"ff0683ff",
   422 => x"e0800c52",
   423 => x"52028c05",
   424 => x"0d0402f8",
   425 => x"050d7370",
   426 => x"902b7190",
   427 => x"2a0783ff",
   428 => x"e0800c52",
   429 => x"0288050d",
   430 => x"0402f405",
   431 => x"0d747652",
   432 => x"53807125",
   433 => x"90387052",
   434 => x"72708405",
   435 => x"5408ff13",
   436 => x"535171f4",
   437 => x"38028c05",
   438 => x"0d0402dc",
   439 => x"050d7a7c",
   440 => x"5a57810b",
   441 => x"a08095d8",
   442 => x"57558358",
   443 => x"7508770c",
   444 => x"76087608",
   445 => x"55537274",
   446 => x"2e8f3873",
   447 => x"52a08095",
   448 => x"e851a080",
   449 => x"828f2d80",
   450 => x"55785276",
   451 => x"51a0808d",
   452 => x"b92d7608",
   453 => x"5372742e",
   454 => x"8f387352",
   455 => x"a080969c",
   456 => x"51a08082",
   457 => x"8f2d8055",
   458 => x"ff188417",
   459 => x"57587780",
   460 => x"25ffb938",
   461 => x"7483ffe0",
   462 => x"800c02a4",
   463 => x"050d0402",
   464 => x"cc050d7e",
   465 => x"a08096d0",
   466 => x"525ba080",
   467 => x"828f2d80",
   468 => x"e1b3578e",
   469 => x"5c76598f",
   470 => x"ffff5a76",
   471 => x"bfffff06",
   472 => x"77107096",
   473 => x"2a708106",
   474 => x"51575858",
   475 => x"74802e85",
   476 => x"38768107",
   477 => x"5776952a",
   478 => x"70810651",
   479 => x"5574802e",
   480 => x"85387681",
   481 => x"325776bf",
   482 => x"ffff0678",
   483 => x"84291c79",
   484 => x"710c5670",
   485 => x"84291c56",
   486 => x"750c7610",
   487 => x"70962a70",
   488 => x"81065156",
   489 => x"5774802e",
   490 => x"85387681",
   491 => x"07577695",
   492 => x"2a708106",
   493 => x"51557480",
   494 => x"2e853876",
   495 => x"813257ff",
   496 => x"1a5a7980",
   497 => x"25ff9438",
   498 => x"78578fff",
   499 => x"ff5a76bf",
   500 => x"ffff0677",
   501 => x"1070962a",
   502 => x"70810651",
   503 => x"57585974",
   504 => x"802e8538",
   505 => x"76810757",
   506 => x"76952a70",
   507 => x"81065155",
   508 => x"74802e85",
   509 => x"38768132",
   510 => x"5776bfff",
   511 => x"ff067984",
   512 => x"291c7008",
   513 => x"57575874",
   514 => x"792e9438",
   515 => x"80760855",
   516 => x"79547953",
   517 => x"a08096e4",
   518 => x"525da080",
   519 => x"828f2d77",
   520 => x"84291b70",
   521 => x"08565674",
   522 => x"782e9438",
   523 => x"80760855",
   524 => x"78547853",
   525 => x"a08096e4",
   526 => x"525da080",
   527 => x"828f2d76",
   528 => x"1070962a",
   529 => x"70810651",
   530 => x"56577480",
   531 => x"2e853876",
   532 => x"81075776",
   533 => x"952a7081",
   534 => x"06515574",
   535 => x"802e8538",
   536 => x"76813257",
   537 => x"ff1a5a79",
   538 => x"8025fee2",
   539 => x"38ff1c5c",
   540 => x"7bfde238",
   541 => x"7c83ffe0",
   542 => x"800c02b4",
   543 => x"050d0402",
   544 => x"cc050d7e",
   545 => x"5b815c80",
   546 => x"5a80c07c",
   547 => x"585d85aa",
   548 => x"d6d5aa7b",
   549 => x"0c7b5881",
   550 => x"56975576",
   551 => x"7607822b",
   552 => x"7b115154",
   553 => x"85aad6d5",
   554 => x"aa740c75",
   555 => x"10ff1656",
   556 => x"56748025",
   557 => x"e6387610",
   558 => x"81195957",
   559 => x"987825d7",
   560 => x"387f527a",
   561 => x"51a0808d",
   562 => x"b92d8157",
   563 => x"ff87c3e1",
   564 => x"f07b0c97",
   565 => x"58807782",
   566 => x"2b7c1170",
   567 => x"0857575a",
   568 => x"5673ff87",
   569 => x"c3e1f02e",
   570 => x"0981068c",
   571 => x"38757a78",
   572 => x"075b5ca0",
   573 => x"80929504",
   574 => x"74085473",
   575 => x"85aad6d5",
   576 => x"aa2e9238",
   577 => x"75750854",
   578 => x"7953a080",
   579 => x"9788525c",
   580 => x"a080828f",
   581 => x"2d7610ff",
   582 => x"19595777",
   583 => x"8025ffb5",
   584 => x"3879802e",
   585 => x"9e387982",
   586 => x"2b52a080",
   587 => x"97a451a0",
   588 => x"80828f2d",
   589 => x"791087ff",
   590 => x"fffe067d",
   591 => x"812c5e5a",
   592 => x"79f2387c",
   593 => x"52a08097",
   594 => x"bc51a080",
   595 => x"828f2d7b",
   596 => x"83ffe080",
   597 => x"0c02b405",
   598 => x"0d0402f8",
   599 => x"050d88bd",
   600 => x"0bff880c",
   601 => x"a0805280",
   602 => x"51a0808d",
   603 => x"da2d83ff",
   604 => x"e0800880",
   605 => x"2e8b38a0",
   606 => x"8097f851",
   607 => x"a080828f",
   608 => x"2da08052",
   609 => x"8051a080",
   610 => x"90ff2d83",
   611 => x"ffe08008",
   612 => x"802e8b38",
   613 => x"a080989c",
   614 => x"51a08082",
   615 => x"8f2d8051",
   616 => x"a0808ebf",
   617 => x"2d83ffe0",
   618 => x"8008802e",
   619 => x"8b38a080",
   620 => x"98b451a0",
   621 => x"80828f2d",
   622 => x"800b83ff",
   623 => x"e0800c02",
   624 => x"88050d04",
   625 => x"00ffffff",
   626 => x"ff00ffff",
   627 => x"ffff00ff",
   628 => x"ffffff00",
   629 => x"30313233",
   630 => x"34353637",
   631 => x"38394142",
   632 => x"43444546",
   633 => x"00000000",
   634 => x"53444843",
   635 => x"20496e69",
   636 => x"7469616c",
   637 => x"697a6174",
   638 => x"696f6e20",
   639 => x"6572726f",
   640 => x"72210a00",
   641 => x"434d4435",
   642 => x"38202564",
   643 => x"0a202000",
   644 => x"434d4435",
   645 => x"385f3220",
   646 => x"25640a20",
   647 => x"20000000",
   648 => x"44657465",
   649 => x"726d696e",
   650 => x"65642053",
   651 => x"44484320",
   652 => x"73746174",
   653 => x"75730a00",
   654 => x"53656e74",
   655 => x"20726573",
   656 => x"65742063",
   657 => x"6f6d6d61",
   658 => x"6e640a00",
   659 => x"53442063",
   660 => x"61726420",
   661 => x"696e6974",
   662 => x"69616c69",
   663 => x"7a617469",
   664 => x"6f6e2065",
   665 => x"72726f72",
   666 => x"210a0000",
   667 => x"43617264",
   668 => x"20726573",
   669 => x"706f6e64",
   670 => x"65642074",
   671 => x"6f207265",
   672 => x"7365740a",
   673 => x"00000000",
   674 => x"53444843",
   675 => x"20636172",
   676 => x"64206465",
   677 => x"74656374",
   678 => x"65640a00",
   679 => x"53656e64",
   680 => x"696e6720",
   681 => x"636d6431",
   682 => x"360a0000",
   683 => x"496e6974",
   684 => x"20646f6e",
   685 => x"650a0000",
   686 => x"52656164",
   687 => x"20636f6d",
   688 => x"6d616e64",
   689 => x"20666169",
   690 => x"6c656420",
   691 => x"61742025",
   692 => x"64202825",
   693 => x"64290a00",
   694 => x"00000000",
   695 => x"55555555",
   696 => x"aaaaaaaa",
   697 => x"ffffffff",
   698 => x"53616e69",
   699 => x"74792063",
   700 => x"6865636b",
   701 => x"20666169",
   702 => x"6c656420",
   703 => x"28626566",
   704 => x"6f726520",
   705 => x"63616368",
   706 => x"65207265",
   707 => x"66726573",
   708 => x"6829206f",
   709 => x"6e202564",
   710 => x"0a000000",
   711 => x"53616e69",
   712 => x"74792063",
   713 => x"6865636b",
   714 => x"20666169",
   715 => x"6c656420",
   716 => x"28616674",
   717 => x"65722063",
   718 => x"61636865",
   719 => x"20726566",
   720 => x"72657368",
   721 => x"29206f6e",
   722 => x"2025640a",
   723 => x"00000000",
   724 => x"43686563",
   725 => x"6b696e67",
   726 => x"206d656d",
   727 => x"6f72792e",
   728 => x"2e2e0a00",
   729 => x"4572726f",
   730 => x"72206174",
   731 => x"2025642c",
   732 => x"20657870",
   733 => x"65637465",
   734 => x"64202564",
   735 => x"2c20676f",
   736 => x"74202564",
   737 => x"0a000000",
   738 => x"42616420",
   739 => x"64617461",
   740 => x"20666f75",
   741 => x"6e642061",
   742 => x"74202564",
   743 => x"20282564",
   744 => x"290a0000",
   745 => x"416c6961",
   746 => x"73657320",
   747 => x"666f756e",
   748 => x"64206174",
   749 => x"2025640a",
   750 => x"00000000",
   751 => x"53445241",
   752 => x"4d207369",
   753 => x"7a652028",
   754 => x"61737375",
   755 => x"6d696e67",
   756 => x"206e6f20",
   757 => x"61646472",
   758 => x"65737320",
   759 => x"6661756c",
   760 => x"74732920",
   761 => x"69732025",
   762 => x"64206d65",
   763 => x"67616279",
   764 => x"7465730a",
   765 => x"00000000",
   766 => x"46697273",
   767 => x"74207374",
   768 => x"61676520",
   769 => x"73616e69",
   770 => x"74792063",
   771 => x"6865636b",
   772 => x"20706173",
   773 => x"7365642e",
   774 => x"0a000000",
   775 => x"41646472",
   776 => x"65737320",
   777 => x"63686563",
   778 => x"6b207061",
   779 => x"73736564",
   780 => x"2e0a0000",
   781 => x"4c465352",
   782 => x"20636865",
   783 => x"636b2070",
   784 => x"61737365",
   785 => x"642e0a00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

